`ifndef COEFFICIENTS_FX_SV_
`define COEFFICIENTS_FX_SV_

package Coefficients_Fx;

	localparam N = 4;
	localparam M = 4;
	localparam COEFF_BIAS = 48;
	localparam logic signed[63:0] Lfr[0:3] = {64'd279328808984837, 64'd279328808984837, 64'd276620165905596, 64'd276620165905596};

	localparam logic signed[63:0] Lfi[0:3] = {64'd9678520698973, - 64'd9678520698973, 64'd3897284466146, - 64'd3897284466146};

	localparam logic signed[63:0] Lbr[0:3] = {64'd279328808984837, 64'd279328808984837, 64'd276620165905596, 64'd276620165905596};

	localparam logic signed[63:0] Lbi[0:3] = {64'd9678520698973, - 64'd9678520698973, 64'd3897284466146, - 64'd3897284466146};

	localparam logic signed[63:0] Wfr[0:3] = {- 64'd969817770, - 64'd969817770, 64'd288523161, 64'd288523161};

	localparam logic signed[63:0] Wfi[0:3] = {- 64'd37246664, 64'd37246664, 64'd555624089, - 64'd555624089};

	localparam logic signed[63:0] Wbr[0:3] = {64'd969817770, 64'd969817770, - 64'd288523161, - 64'd288523161};

	localparam logic signed[63:0] Wbi[0:3] = {64'd37246664, - 64'd37246664, - 64'd555624089, 64'd555624089};

	localparam logic signed[63:0] Ffr[0:3][0:79] = '{
		'{- 64'd140566688200280032, - 64'd9885414325770184, 64'd784783703179973, - 64'd5825088699075, - 64'd145386281648678336, - 64'd9392113046470502, 64'd788209301998607, - 64'd7194786936037, - 64'd149958010880262208, - 64'd8894071819875330, 64'd790609165282370, - 64'd8536372222145, - 64'd154279677146064768, - 64'd8391974850718128, 64'd791994685585595, - 64'd9848574200773, - 64'd158349422693806176, - 64'd7886501789734974, 64'd792378354122056, - 64'd11130176760670, - 64'd162165728295357504, - 64'd7378326954378150, 64'd791773729878953, - 64'd12380018784571, - 64'd165727410388915104, - 64'd6868118567062459, 64'd790195407839052, - 64'd13596994819126, - 64'd169033617844827264, - 64'd6356538011643610, 64'd787658986362872, - 64'd14780055666371, - 64'd172083828364358208, - 64'd5844239108795604, 64'd784181033783172, - 64'd15928208897149, - 64'd174877844520997888, - 64'd5331867410921166, 64'd779779054264189, - 64'd17040519286910, - 64'd177415789454236576, - 64'd4820059517196292, 64'd774471452978286, - 64'd18116109174444, - 64'd179698102226013728, - 64'd4309442409316473, 64'd768277500652777, - 64'd19154158744190, - 64'd181725532850327872, - 64'd3800632808478583, 64'd761217297539715, - 64'd20153906232826, - 64'd183499137006750880, - 64'd3294236554098600, 64'd753311736861436, - 64'd21114648060965, - 64'd185020270448833216, - 64'd2790848004731313, 64'd744582467784540, - 64'd22035738890815, - 64'd186290583118609664, - 64'd2291049461624139, 64'd735051857974838, - 64'd22916591610800, - 64'd187312012978625216, - 64'd1795410615303047, 64'd724742955785610, - 64'd23756677248161, - 64'd188086779573087232, - 64'd1304488015554396, 64'd713679452131176, - 64'd24555524810658, - 64'd188617377329927840, - 64'd818824565132426, 64'd701885642097519, - 64'd25312721058582, - 64'd188906568615713280, - 64'd338949037488046, 64'd689386386341246, - 64'd26027910208299},
		'{- 64'd140566688200270224, - 64'd9885414325770250, 64'd784783703180054, - 64'd5825088699114, - 64'd145386281648669024, - 64'd9392113046470558, 64'd788209301998685, - 64'd7194786936074, - 64'd149958010880253376, - 64'd8894071819875381, 64'd790609165282444, - 64'd8536372222180, - 64'd154279677146056416, - 64'd8391974850718170, 64'd791994685585666, - 64'd9848574200808, - 64'd158349422693798304, - 64'd7886501789735009, 64'd792378354122124, - 64'd11130176760702, - 64'd162165728295350112, - 64'd7378326954378176, 64'd791773729879019, - 64'd12380018784603, - 64'd165727410388908224, - 64'd6868118567062478, 64'd790195407839114, - 64'd13596994819156, - 64'd169033617844820864, - 64'd6356538011643622, 64'd787658986362931, - 64'd14780055666399, - 64'd172083828364352320, - 64'd5844239108795608, 64'd784181033783228, - 64'd15928208897176, - 64'd174877844520992512, - 64'd5331867410921162, 64'd779779054264242, - 64'd17040519286936, - 64'd177415789454231680, - 64'd4820059517196282, 64'd774471452978336, - 64'd18116109174468, - 64'd179698102226009312, - 64'd4309442409316455, 64'd768277500652824, - 64'd19154158744212, - 64'd181725532850323968, - 64'd3800632808478558, 64'd761217297539758, - 64'd20153906232847, - 64'd183499137006747456, - 64'd3294236554098568, 64'd753311736861476, - 64'd21114648060984, - 64'd185020270448830272, - 64'd2790848004731274, 64'd744582467784576, - 64'd22035738890833, - 64'd186290583118607232, - 64'd2291049461624093, 64'd735051857974872, - 64'd22916591610817, - 64'd187312012978623264, - 64'd1795410615302995, 64'd724742955785640, - 64'd23756677248175, - 64'd188086779573085760, - 64'd1304488015554337, 64'd713679452131203, - 64'd24555524810672, - 64'd188617377329926816, - 64'd818824565132361, 64'd701885642097543, - 64'd25312721058593, - 64'd188906568615712736, - 64'd338949037487975, 64'd689386386341266, - 64'd26027910208309},
		'{64'd140075906892424448, 64'd9853761721326258, - 64'd764775131297287, 64'd74640218037739, 64'd144883670460580832, 64'd9379232192999704, - 64'd734786646196608, 64'd72645337313765, 64'd149457063372826912, 64'd8916251390512551, - 64'd705458504944230, 64'd70682757393738, 64'd153801818429928864, 64'd8464653072160863, - 64'd676782598859692, 64'd68752339930603, 64'd157923585329725408, 64'd8024271081254372, - 64'd648750775938709, 64'd66853935548267, 64'd161827930729348224, 64'd7594939424508485, - 64'd621354846314382, 64'd64987384289729, 64'd165520338345949696, 64'd7176492347690528, - 64'd594586587551199, 64'd63152516055151, 64'd169006209094579136, 64'd6768764408576604, - 64'd568437749774955, 64'd61349151029988, 64'd172290861261876608, 64'd6371590547274816, - 64'd542900060641629, 64'd59577100103315, 64'd175379530714281344, 64'd5984806153970032, - 64'd517965230148294, 64'd57836165276473, 64'd178277371139479776, 64'd5608247134144710, - 64'd493624955289057, 64'd56126140062170, 64'd180989454319843648, 64'd5241749971329742, - 64'd469870924559030, 64'd54446809874161, 64'd183520770436637568, 64'd4885151787438578, - 64'd446694822309294, 64'd52797952407633, 64'd185876228403800256, 64'd4538290400737318, - 64'd424088332955797, 64'd51179338010443, 64'd188060656230130816, 64'd4201004381502817, - 64'd402043145045090, 64'd49590730045313, 64'd190078801408736576, 64'd3873133105420170, - 64'd380550955179780, 64'd48031885243131, 64'd191935331332625312, 64'd3554516804770342, - 64'd359603471806553, 64'd46502554047483, 64'd193634833735349216, 64'd3244996617458062, - 64'd339192418869587, 64'd45002480950541, 64'd195181817155633024, 64'd2944414633929432, - 64'd319309539332144, 64'd43531404820443, 64'd196580711424943872, 64'd2652613942028054, - 64'd299946598569100, 64'd42089059220290},
		'{64'd140075906892391456, 64'd9853761721326572, - 64'd764775131297532, 64'd74640218037855, 64'd144883670460548576, 64'd9379232193000008, - 64'd734786646196848, 64'd72645337313879, 64'd149457063372795392, 64'd8916251390512847, - 64'd705458504944465, 64'd70682757393850, 64'd153801818429898048, 64'd8464653072161152, - 64'd676782598859921, 64'd68752339930712, 64'd157923585329695264, 64'd8024271081254654, - 64'd648750775938934, 64'd66853935548374, 64'd161827930729318784, 64'd7594939424508759, - 64'd621354846314602, 64'd64987384289833, 64'd165520338345920960, 64'd7176492347690794, - 64'd594586587551414, 64'd63152516055253, 64'd169006209094551104, 64'd6768764408576861, - 64'd568437749775165, 64'd61349151030088, 64'd172290861261849184, 64'd6371590547275066, - 64'd542900060641834, 64'd59577100103412, 64'd175379530714254592, 64'd5984806153970275, - 64'd517965230148495, 64'd57836165276568, 64'd178277371139453696, 64'd5608247134144946, - 64'd493624955289254, 64'd56126140062264, 64'd180989454319818176, 64'd5241749971329970, - 64'd469870924559222, 64'd54446809874252, 64'd183520770436612736, 64'd4885151787438800, - 64'd446694822309481, 64'd52797952407722, 64'd185876228403776064, 64'd4538290400737533, - 64'd424088332955980, 64'd51179338010530, 64'd188060656230107200, 64'd4201004381503025, - 64'd402043145045268, 64'd49590730045398, 64'd190078801408713600, 64'd3873133105420372, - 64'd380550955179954, 64'd48031885243214, 64'd191935331332602912, 64'd3554516804770536, - 64'd359603471806723, 64'd46502554047563, 64'd193634833735327424, 64'd3244996617458250, - 64'd339192418869753, 64'd45002480950620, 64'd195181817155611776, 64'd2944414633929615, - 64'd319309539332306, 64'd43531404820520, 64'd196580711424923200, 64'd2652613942028230, - 64'd299946598569257, 64'd42089059220365}};

	localparam logic signed[63:0] Ffi[0:3][0:79] = '{
		'{64'd171335547524263200, - 64'd12154358354823768, - 64'd273646963785454, 64'd41125850643455, 64'd165195774660932896, - 64'd12401594881331294, - 64'd244575684721808, 64'd40611981820778, 64'd158937094060300544, - 64'd12629984127848390, - 64'd215608276745190, 64'd40054934012185, 64'd152568935174788992, - 64'd12839506816448324, - 64'd186779217797280, 64'd39456003109506, 64'd146100731163903456, - 64'd13030167342581730, - 64'd158122331201997, 64'd38816518804988, 64'd139541907140790608, - 64'd13201993437984464, - 64'd129670752879361, 64'd38137842468350, 64'd132901868593432608, - 64'd13355035809359964, - 64'd101456899871346, 64'd37421365014280, 64'd126189989992392256, - 64'd13489367753623618, - 64'd73512440200407, 64'd36668504763159, 64'd119415603596628576, - 64'd13605084750514794, - 64'd45868264079387, 64'd35880705297761, 64'd112587988468493120, - 64'd13702304033398926, - 64'd18554456489584, 64'd35059433318633, 64'd105716359708603408, - 64'd13781164139097620, 64'd8399728858155, 64'd34206176500850, 64'd98809857920867184, - 64'd13841824437598938, 64'd34965894166412, 64'd33322441354776, 64'd91877538917501568, - 64'd13884464642513178, 64'd61116520787212, 64'd32409751093424, 64'd84928363673455136, - 64'd13909284303151072, 64'd86824991041977, 64'd31469643508976, 64'd77971188539201072, - 64'd13916502279111976, 64'd112065608618179, 64'd30503668860966, 64'd71014755720421544, - 64'd13906356198278744, 64'd136813617537335, 64'd29513387778584, 64'd64067684032655120, - 64'd13879101899124208, 64'd161045219690830, 64'd28500369179499, 64'd57138459938522864, - 64'd13835012858240672, 64'd184737590941875, 64'd27466188207556, 64'd50235428874693296, - 64'd13774379604009744, 64'd207868895793713, 64'd26412424191648, 64'd43366786875285072, - 64'd13697509117333812, 64'd230418300625970, 64'd25340658627977},
		'{- 64'd171335547524274880, 64'd12154358354823986, 64'd273646963785388, - 64'd41125850643424, - 64'd165195774660944832, 64'd12401594881331512, 64'd244575684721740, - 64'd40611981820746, - 64'd158937094060312704, 64'd12629984127848608, 64'd215608276745120, - 64'd40054934012152, - 64'd152568935174801344, 64'd12839506816448544, 64'd186779217797207, - 64'd39456003109472, - 64'd146100731163916000, 64'd13030167342581948, 64'd158122331201923, - 64'd38816518804953, - 64'd139541907140803344, 64'd13201993437984680, 64'd129670752879284, - 64'd38137842468314, - 64'd132901868593445488, 64'd13355035809360184, 64'd101456899871268, - 64'd37421365014244, - 64'd126189989992405280, 64'd13489367753623834, 64'd73512440200328, - 64'd36668504763122, - 64'd119415603596641744, 64'd13605084750515008, 64'd45868264079306, - 64'd35880705297723, - 64'd112587988468506368, 64'd13702304033399140, 64'd18554456489502, - 64'd35059433318594, - 64'd105716359708616752, 64'd13781164139097830, - 64'd8399728858238, - 64'd34206176500811, - 64'd98809857920880608, 64'd13841824437599146, - 64'd34965894166496, - 64'd33322441354737, - 64'd91877538917515024, 64'd13884464642513384, - 64'd61116520787298, - 64'd32409751093384, - 64'd84928363673468624, 64'd13909284303151278, - 64'd86824991042064, - 64'd31469643508935, - 64'd77971188539214592, 64'd13916502279112180, - 64'd112065608618266, - 64'd30503668860925, - 64'd71014755720435040, 64'd13906356198278946, - 64'd136813617537422, - 64'd29513387778543, - 64'd64067684032668600, 64'd13879101899124402, - 64'd161045219690918, - 64'd28500369179458, - 64'd57138459938536304, 64'd13835012858240864, - 64'd184737590941963, - 64'd27466188207515, - 64'd50235428874706688, 64'd13774379604009932, - 64'd207868895793802, - 64'd26412424191606, - 64'd43366786875298400, 64'd13697509117334000, - 64'd230418300626059, - 64'd25340658627935},
		'{- 64'd521724083101841984, 64'd21997377867528308, - 64'd1213195910000991, 64'd51098366062182, - 64'd510786033091518720, 64'd21754407085315836, - 64'd1202860034296424, 64'd51250497747666, - 64'd499970071877531520, 64'd21509056697681584, - 64'd1192287210580083, 64'd51372384512954, - 64'd489277338783569856, 64'd21261527650388452, - 64'd1181490668751241, 64'd51464995249811, - 64'd478708874106558464, 64'd21012015121564524, - 64'd1170483298250872, 64'd51529280223250, - 64'd468265621975284032, 64'd20760708622358940, - 64'd1159277653333931, 64'd51566171240098, - 64'd457948433158855872, 64'd20507792096947004, - 64'd1147885958326313, 64'd51576581820854, - 64'd447758067825332544, 64'd20253444021857912, - 64'd1136320112864451, 64'd51561407374649, - 64'd437695198250858304, 64'd19997837504599376, - 64'd1124591697115560, 64'd51521525377118, - 64'd427760411479669376, 64'd19741140381554972, - 64'd1112711976976651, 64'd51457795550997, - 64'd417954211935337216, 64'd19483515315130860, - 64'd1100691909250479, 64'd51371060049257, - 64'd408277023983631488, 64'd19225119890130096, - 64'd1088542146796688, 64'd51262143640617, - 64'd398729194447392384, 64'd18966106709333468, - 64'd1076273043656470, 64'd51131853897238, - 64'd389310995073816128, 64'd18706623488267196, - 64'd1063894660149130, 64'd50980981384460, - 64'd380022624954562880, 64'd18446813149138748, - 64'd1051416767939034, 64'd50810299852398, - 64'd370864212899109312, 64'd18186813913923108, - 64'd1038848855071444, 64'd50620566429252, - 64'd361835819761773056, 64'd17926759396582846, - 64'd1026200130975855, 64'd50412521816173, - 64'd352937440722847296, 64'd17666778694406360, - 64'd1013479531435485, 64'd50186890483540, - 64'd344169007524289984, 64'd17406996478449558, - 64'd1000695723521634, 64'd49944380868501, - 64'd335530390660419200, 64'd17147533083067242, - 64'd987857110491698, 64'd49685685573640},
		'{64'd521724083101853696, - 64'd21997377867528528, 64'd1213195910001057, - 64'd51098366062212, 64'd510786033091530688, - 64'd21754407085316056, 64'd1202860034296492, - 64'd51250497747698, 64'd499970071877543744, - 64'd21509056697681804, 64'd1192287210580153, - 64'd51372384512987, 64'd489277338783582272, - 64'd21261527650388672, 64'd1181490668751314, - 64'd51464995249844, 64'd478708874106571072, - 64'd21012015121564748, 64'd1170483298250947, - 64'd51529280223284, 64'd468265621975296832, - 64'd20760708622359164, 64'd1159277653334007, - 64'd51566171240133, 64'd457948433158868928, - 64'd20507792096947228, 64'd1147885958326391, - 64'd51576581820890, 64'd447758067825345728, - 64'd20253444021858132, 64'd1136320112864531, - 64'd51561407374686, 64'd437695198250871680, - 64'd19997837504599600, 64'd1124591697115642, - 64'd51521525377156, 64'd427760411479682880, - 64'd19741140381555192, 64'd1112711976976734, - 64'd51457795551035, 64'd417954211935350912, - 64'd19483515315131080, 64'd1100691909250563, - 64'd51371060049297, 64'd408277023983645248, - 64'd19225119890130312, 64'd1088542146796774, - 64'd51262143640657, 64'd398729194447406272, - 64'd18966106709333684, 64'd1076273043656556, - 64'd51131853897278, 64'd389310995073830080, - 64'd18706623488267416, 64'd1063894660149218, - 64'd50980981384501, 64'd380022624954576960, - 64'd18446813149138968, 64'd1051416767939123, - 64'd50810299852440, 64'd370864212899123520, - 64'd18186813913923328, 64'd1038848855071534, - 64'd50620566429294, 64'd361835819761787264, - 64'd17926759396583062, 64'd1026200130975946, - 64'd50412521816215, 64'd352937440722861568, - 64'd17666778694406576, 64'd1013479531435576, - 64'd50186890483582, 64'd344169007524304384, - 64'd17406996478449772, 64'd1000695723521726, - 64'd49944380868544, 64'd335530390660433600, - 64'd17147533083067456, 64'd987857110491791, - 64'd49685685573683}};

	localparam logic signed[63:0] Fbr[0:3][0:79] = '{
		'{64'd140566688200280032, - 64'd9885414325770184, - 64'd784783703179973, - 64'd5825088699075, 64'd145386281648678336, - 64'd9392113046470502, - 64'd788209301998607, - 64'd7194786936037, 64'd149958010880262208, - 64'd8894071819875330, - 64'd790609165282370, - 64'd8536372222145, 64'd154279677146064768, - 64'd8391974850718128, - 64'd791994685585595, - 64'd9848574200773, 64'd158349422693806176, - 64'd7886501789734974, - 64'd792378354122056, - 64'd11130176760670, 64'd162165728295357504, - 64'd7378326954378150, - 64'd791773729878953, - 64'd12380018784571, 64'd165727410388915104, - 64'd6868118567062459, - 64'd790195407839052, - 64'd13596994819126, 64'd169033617844827264, - 64'd6356538011643610, - 64'd787658986362872, - 64'd14780055666371, 64'd172083828364358208, - 64'd5844239108795604, - 64'd784181033783172, - 64'd15928208897149, 64'd174877844520997888, - 64'd5331867410921166, - 64'd779779054264189, - 64'd17040519286910, 64'd177415789454236576, - 64'd4820059517196292, - 64'd774471452978286, - 64'd18116109174444, 64'd179698102226013728, - 64'd4309442409316473, - 64'd768277500652777, - 64'd19154158744190, 64'd181725532850327872, - 64'd3800632808478583, - 64'd761217297539715, - 64'd20153906232826, 64'd183499137006750880, - 64'd3294236554098600, - 64'd753311736861436, - 64'd21114648060965, 64'd185020270448833216, - 64'd2790848004731313, - 64'd744582467784540, - 64'd22035738890815, 64'd186290583118609664, - 64'd2291049461624139, - 64'd735051857974838, - 64'd22916591610800, 64'd187312012978625216, - 64'd1795410615303047, - 64'd724742955785610, - 64'd23756677248161, 64'd188086779573087232, - 64'd1304488015554396, - 64'd713679452131176, - 64'd24555524810658, 64'd188617377329927840, - 64'd818824565132426, - 64'd701885642097519, - 64'd25312721058582, 64'd188906568615713280, - 64'd338949037488046, - 64'd689386386341246, - 64'd26027910208299},
		'{64'd140566688200270224, - 64'd9885414325770250, - 64'd784783703180054, - 64'd5825088699114, 64'd145386281648669024, - 64'd9392113046470558, - 64'd788209301998685, - 64'd7194786936074, 64'd149958010880253376, - 64'd8894071819875381, - 64'd790609165282444, - 64'd8536372222180, 64'd154279677146056416, - 64'd8391974850718170, - 64'd791994685585666, - 64'd9848574200808, 64'd158349422693798304, - 64'd7886501789735009, - 64'd792378354122124, - 64'd11130176760702, 64'd162165728295350112, - 64'd7378326954378176, - 64'd791773729879019, - 64'd12380018784603, 64'd165727410388908224, - 64'd6868118567062478, - 64'd790195407839114, - 64'd13596994819156, 64'd169033617844820864, - 64'd6356538011643622, - 64'd787658986362931, - 64'd14780055666399, 64'd172083828364352320, - 64'd5844239108795608, - 64'd784181033783228, - 64'd15928208897176, 64'd174877844520992512, - 64'd5331867410921162, - 64'd779779054264242, - 64'd17040519286936, 64'd177415789454231680, - 64'd4820059517196282, - 64'd774471452978336, - 64'd18116109174468, 64'd179698102226009312, - 64'd4309442409316455, - 64'd768277500652824, - 64'd19154158744212, 64'd181725532850323968, - 64'd3800632808478558, - 64'd761217297539758, - 64'd20153906232847, 64'd183499137006747456, - 64'd3294236554098568, - 64'd753311736861476, - 64'd21114648060984, 64'd185020270448830272, - 64'd2790848004731274, - 64'd744582467784576, - 64'd22035738890833, 64'd186290583118607232, - 64'd2291049461624093, - 64'd735051857974872, - 64'd22916591610817, 64'd187312012978623264, - 64'd1795410615302995, - 64'd724742955785640, - 64'd23756677248175, 64'd188086779573085760, - 64'd1304488015554337, - 64'd713679452131203, - 64'd24555524810672, 64'd188617377329926816, - 64'd818824565132361, - 64'd701885642097543, - 64'd25312721058593, 64'd188906568615712736, - 64'd338949037487975, - 64'd689386386341266, - 64'd26027910208309},
		'{- 64'd140075906892424448, 64'd9853761721326258, 64'd764775131297287, 64'd74640218037739, - 64'd144883670460580832, 64'd9379232192999704, 64'd734786646196608, 64'd72645337313765, - 64'd149457063372826912, 64'd8916251390512551, 64'd705458504944230, 64'd70682757393738, - 64'd153801818429928864, 64'd8464653072160863, 64'd676782598859692, 64'd68752339930603, - 64'd157923585329725408, 64'd8024271081254372, 64'd648750775938709, 64'd66853935548267, - 64'd161827930729348224, 64'd7594939424508485, 64'd621354846314382, 64'd64987384289729, - 64'd165520338345949696, 64'd7176492347690528, 64'd594586587551199, 64'd63152516055151, - 64'd169006209094579136, 64'd6768764408576604, 64'd568437749774955, 64'd61349151029988, - 64'd172290861261876608, 64'd6371590547274816, 64'd542900060641629, 64'd59577100103315, - 64'd175379530714281344, 64'd5984806153970032, 64'd517965230148294, 64'd57836165276473, - 64'd178277371139479776, 64'd5608247134144710, 64'd493624955289057, 64'd56126140062170, - 64'd180989454319843648, 64'd5241749971329742, 64'd469870924559030, 64'd54446809874161, - 64'd183520770436637568, 64'd4885151787438578, 64'd446694822309294, 64'd52797952407633, - 64'd185876228403800256, 64'd4538290400737318, 64'd424088332955797, 64'd51179338010443, - 64'd188060656230130816, 64'd4201004381502817, 64'd402043145045090, 64'd49590730045313, - 64'd190078801408736576, 64'd3873133105420170, 64'd380550955179780, 64'd48031885243131, - 64'd191935331332625312, 64'd3554516804770342, 64'd359603471806553, 64'd46502554047483, - 64'd193634833735349216, 64'd3244996617458062, 64'd339192418869587, 64'd45002480950541, - 64'd195181817155633024, 64'd2944414633929432, 64'd319309539332144, 64'd43531404820443, - 64'd196580711424943872, 64'd2652613942028054, 64'd299946598569100, 64'd42089059220290},
		'{- 64'd140075906892391456, 64'd9853761721326572, 64'd764775131297532, 64'd74640218037855, - 64'd144883670460548576, 64'd9379232193000008, 64'd734786646196848, 64'd72645337313879, - 64'd149457063372795392, 64'd8916251390512847, 64'd705458504944465, 64'd70682757393850, - 64'd153801818429898048, 64'd8464653072161152, 64'd676782598859921, 64'd68752339930712, - 64'd157923585329695264, 64'd8024271081254654, 64'd648750775938934, 64'd66853935548374, - 64'd161827930729318784, 64'd7594939424508759, 64'd621354846314602, 64'd64987384289833, - 64'd165520338345920960, 64'd7176492347690794, 64'd594586587551414, 64'd63152516055253, - 64'd169006209094551104, 64'd6768764408576861, 64'd568437749775165, 64'd61349151030088, - 64'd172290861261849184, 64'd6371590547275066, 64'd542900060641834, 64'd59577100103412, - 64'd175379530714254592, 64'd5984806153970275, 64'd517965230148495, 64'd57836165276568, - 64'd178277371139453696, 64'd5608247134144946, 64'd493624955289254, 64'd56126140062264, - 64'd180989454319818176, 64'd5241749971329970, 64'd469870924559222, 64'd54446809874252, - 64'd183520770436612736, 64'd4885151787438800, 64'd446694822309481, 64'd52797952407722, - 64'd185876228403776064, 64'd4538290400737533, 64'd424088332955980, 64'd51179338010530, - 64'd188060656230107200, 64'd4201004381503025, 64'd402043145045268, 64'd49590730045398, - 64'd190078801408713600, 64'd3873133105420372, 64'd380550955179954, 64'd48031885243214, - 64'd191935331332602912, 64'd3554516804770536, 64'd359603471806723, 64'd46502554047563, - 64'd193634833735327424, 64'd3244996617458250, 64'd339192418869753, 64'd45002480950620, - 64'd195181817155611776, 64'd2944414633929615, 64'd319309539332306, 64'd43531404820520, - 64'd196580711424923200, 64'd2652613942028230, 64'd299946598569257, 64'd42089059220365}};

	localparam logic signed[63:0] Fbi[0:3][0:79] = '{
		'{- 64'd171335547524263200, - 64'd12154358354823768, 64'd273646963785454, 64'd41125850643455, - 64'd165195774660932896, - 64'd12401594881331294, 64'd244575684721808, 64'd40611981820778, - 64'd158937094060300544, - 64'd12629984127848390, 64'd215608276745190, 64'd40054934012185, - 64'd152568935174788992, - 64'd12839506816448324, 64'd186779217797280, 64'd39456003109506, - 64'd146100731163903456, - 64'd13030167342581730, 64'd158122331201997, 64'd38816518804988, - 64'd139541907140790608, - 64'd13201993437984464, 64'd129670752879361, 64'd38137842468350, - 64'd132901868593432608, - 64'd13355035809359964, 64'd101456899871346, 64'd37421365014280, - 64'd126189989992392256, - 64'd13489367753623618, 64'd73512440200407, 64'd36668504763159, - 64'd119415603596628576, - 64'd13605084750514794, 64'd45868264079387, 64'd35880705297761, - 64'd112587988468493120, - 64'd13702304033398926, 64'd18554456489584, 64'd35059433318633, - 64'd105716359708603408, - 64'd13781164139097620, - 64'd8399728858155, 64'd34206176500850, - 64'd98809857920867184, - 64'd13841824437598938, - 64'd34965894166412, 64'd33322441354776, - 64'd91877538917501568, - 64'd13884464642513178, - 64'd61116520787212, 64'd32409751093424, - 64'd84928363673455136, - 64'd13909284303151072, - 64'd86824991041977, 64'd31469643508976, - 64'd77971188539201072, - 64'd13916502279111976, - 64'd112065608618179, 64'd30503668860966, - 64'd71014755720421544, - 64'd13906356198278744, - 64'd136813617537335, 64'd29513387778584, - 64'd64067684032655120, - 64'd13879101899124208, - 64'd161045219690830, 64'd28500369179499, - 64'd57138459938522864, - 64'd13835012858240672, - 64'd184737590941875, 64'd27466188207556, - 64'd50235428874693296, - 64'd13774379604009744, - 64'd207868895793713, 64'd26412424191648, - 64'd43366786875285072, - 64'd13697509117333812, - 64'd230418300625970, 64'd25340658627977},
		'{64'd171335547524274880, 64'd12154358354823986, - 64'd273646963785388, - 64'd41125850643424, 64'd165195774660944832, 64'd12401594881331512, - 64'd244575684721740, - 64'd40611981820746, 64'd158937094060312704, 64'd12629984127848608, - 64'd215608276745120, - 64'd40054934012152, 64'd152568935174801344, 64'd12839506816448544, - 64'd186779217797207, - 64'd39456003109472, 64'd146100731163916000, 64'd13030167342581948, - 64'd158122331201923, - 64'd38816518804953, 64'd139541907140803344, 64'd13201993437984680, - 64'd129670752879284, - 64'd38137842468314, 64'd132901868593445488, 64'd13355035809360184, - 64'd101456899871268, - 64'd37421365014244, 64'd126189989992405280, 64'd13489367753623834, - 64'd73512440200328, - 64'd36668504763122, 64'd119415603596641744, 64'd13605084750515008, - 64'd45868264079306, - 64'd35880705297723, 64'd112587988468506368, 64'd13702304033399140, - 64'd18554456489502, - 64'd35059433318594, 64'd105716359708616752, 64'd13781164139097830, 64'd8399728858238, - 64'd34206176500811, 64'd98809857920880608, 64'd13841824437599146, 64'd34965894166496, - 64'd33322441354737, 64'd91877538917515024, 64'd13884464642513384, 64'd61116520787298, - 64'd32409751093384, 64'd84928363673468624, 64'd13909284303151278, 64'd86824991042064, - 64'd31469643508935, 64'd77971188539214592, 64'd13916502279112180, 64'd112065608618266, - 64'd30503668860925, 64'd71014755720435040, 64'd13906356198278946, 64'd136813617537422, - 64'd29513387778543, 64'd64067684032668600, 64'd13879101899124402, 64'd161045219690918, - 64'd28500369179458, 64'd57138459938536304, 64'd13835012858240864, 64'd184737590941963, - 64'd27466188207515, 64'd50235428874706688, 64'd13774379604009932, 64'd207868895793802, - 64'd26412424191606, 64'd43366786875298400, 64'd13697509117334000, 64'd230418300626059, - 64'd25340658627935},
		'{64'd521724083101841984, 64'd21997377867528308, 64'd1213195910000991, 64'd51098366062182, 64'd510786033091518720, 64'd21754407085315836, 64'd1202860034296424, 64'd51250497747666, 64'd499970071877531520, 64'd21509056697681584, 64'd1192287210580083, 64'd51372384512954, 64'd489277338783569856, 64'd21261527650388452, 64'd1181490668751241, 64'd51464995249811, 64'd478708874106558464, 64'd21012015121564524, 64'd1170483298250872, 64'd51529280223250, 64'd468265621975284032, 64'd20760708622358940, 64'd1159277653333931, 64'd51566171240098, 64'd457948433158855872, 64'd20507792096947004, 64'd1147885958326313, 64'd51576581820854, 64'd447758067825332544, 64'd20253444021857912, 64'd1136320112864451, 64'd51561407374649, 64'd437695198250858304, 64'd19997837504599376, 64'd1124591697115560, 64'd51521525377118, 64'd427760411479669376, 64'd19741140381554972, 64'd1112711976976651, 64'd51457795550997, 64'd417954211935337216, 64'd19483515315130860, 64'd1100691909250479, 64'd51371060049257, 64'd408277023983631488, 64'd19225119890130096, 64'd1088542146796688, 64'd51262143640617, 64'd398729194447392384, 64'd18966106709333468, 64'd1076273043656470, 64'd51131853897238, 64'd389310995073816128, 64'd18706623488267196, 64'd1063894660149130, 64'd50980981384460, 64'd380022624954562880, 64'd18446813149138748, 64'd1051416767939034, 64'd50810299852398, 64'd370864212899109312, 64'd18186813913923108, 64'd1038848855071444, 64'd50620566429252, 64'd361835819761773056, 64'd17926759396582846, 64'd1026200130975855, 64'd50412521816173, 64'd352937440722847296, 64'd17666778694406360, 64'd1013479531435485, 64'd50186890483540, 64'd344169007524289984, 64'd17406996478449558, 64'd1000695723521634, 64'd49944380868501, 64'd335530390660419200, 64'd17147533083067242, 64'd987857110491698, 64'd49685685573640},
		'{- 64'd521724083101853696, - 64'd21997377867528528, - 64'd1213195910001057, - 64'd51098366062212, - 64'd510786033091530688, - 64'd21754407085316056, - 64'd1202860034296492, - 64'd51250497747698, - 64'd499970071877543744, - 64'd21509056697681804, - 64'd1192287210580153, - 64'd51372384512987, - 64'd489277338783582272, - 64'd21261527650388672, - 64'd1181490668751314, - 64'd51464995249844, - 64'd478708874106571072, - 64'd21012015121564748, - 64'd1170483298250947, - 64'd51529280223284, - 64'd468265621975296832, - 64'd20760708622359164, - 64'd1159277653334007, - 64'd51566171240133, - 64'd457948433158868928, - 64'd20507792096947228, - 64'd1147885958326391, - 64'd51576581820890, - 64'd447758067825345728, - 64'd20253444021858132, - 64'd1136320112864531, - 64'd51561407374686, - 64'd437695198250871680, - 64'd19997837504599600, - 64'd1124591697115642, - 64'd51521525377156, - 64'd427760411479682880, - 64'd19741140381555192, - 64'd1112711976976734, - 64'd51457795551035, - 64'd417954211935350912, - 64'd19483515315131080, - 64'd1100691909250563, - 64'd51371060049297, - 64'd408277023983645248, - 64'd19225119890130312, - 64'd1088542146796774, - 64'd51262143640657, - 64'd398729194447406272, - 64'd18966106709333684, - 64'd1076273043656556, - 64'd51131853897278, - 64'd389310995073830080, - 64'd18706623488267416, - 64'd1063894660149218, - 64'd50980981384501, - 64'd380022624954576960, - 64'd18446813149138968, - 64'd1051416767939123, - 64'd50810299852440, - 64'd370864212899123520, - 64'd18186813913923328, - 64'd1038848855071534, - 64'd50620566429294, - 64'd361835819761787264, - 64'd17926759396583062, - 64'd1026200130975946, - 64'd50412521816215, - 64'd352937440722861568, - 64'd17666778694406576, - 64'd1013479531435576, - 64'd50186890483582, - 64'd344169007524304384, - 64'd17406996478449772, - 64'd1000695723521726, - 64'd49944380868544, - 64'd335530390660433600, - 64'd17147533083067456, - 64'd987857110491791, - 64'd49685685573683}};

	localparam logic signed[63:0] hf[0:1199] = {64'd3360891076608, - 64'd1740072192, - 64'd2258560256, 64'd2309433, 64'd3359151226880, - 64'd5218416128, - 64'd2253798656, 64'd6921711, 64'd3355673624576, - 64'd8691364864, - 64'd2244285696, 64'd11514461, 64'd3350461415424, - 64'd12155332608, - 64'd2230039808, 64'd16075163, 64'd3343520366592, - 64'd15606747136, - 64'd2211088640, 64'd20591730, 64'd3334857293824, - 64'd19042058240, - 64'd2187467776, 64'd25052516, 64'd3324481372160, - 64'd22457741312, - 64'd2159221248, 64'd29446316, 64'd3312403349504, - 64'd25850302464, - 64'd2126401536, 64'd33762368, 64'd3298635546624, - 64'd29216280576, - 64'd2089067776, 64'd37990368, 64'd3283192119296, - 64'd32552259584, - 64'd2047287168, 64'd42120460, 64'd3266088796160, - 64'd35854868480, - 64'd2001134208, 64'd46143240, 64'd3247343403008, - 64'd39120789504, - 64'd1950690048, 64'd50049756, 64'd3226974814208, - 64'd42346749952, - 64'd1896042368, 64'd53831528, 64'd3205003739136, - 64'd45529546752, - 64'd1837285632, 64'd57480512, 64'd3181452984320, - 64'd48666038272, - 64'd1774520192, 64'd60989140, 64'd3156345880576, - 64'd51753148416, - 64'd1707852160, 64'd64350292, 64'd3129708380160, - 64'd54787874816, - 64'd1637393280, 64'd67557296, 64'd3101567221760, - 64'd57767292928, - 64'd1563260672, 64'd70603936, 64'd3071950979072, - 64'd60688547840, - 64'd1485576448, 64'd73484464, 64'd3040889012224, - 64'd63548878848, - 64'd1404467200, 64'd76193552, 64'd3008412516352, - 64'd66345603072, - 64'd1320064256, 64'd78726344, 64'd2974554259456, - 64'd69076131840, - 64'd1232503040, 64'd81078400, 64'd2939347795968, - 64'd71737966592, - 64'd1141922688, 64'd83245736, 64'd2902828253184, - 64'd74328702976, - 64'd1048465984, 64'd85224800, 64'd2865031544832, - 64'd76846030848, - 64'd952279104, 64'd87012456, 64'd2825994895360, - 64'd79287738368, - 64'd853511232, 64'd88605992, 64'd2785756577792, - 64'd81651720192, - 64'd752314240, 64'd90003120, 64'd2744356438016, - 64'd83935985664, - 64'd648842368, 64'd91201968, 64'd2701834321920, - 64'd86138626048, - 64'd543252352, 64'd92201048, 64'd2658231648256, - 64'd88257855488, - 64'd435702464, 64'd92999280, 64'd2613590622208, - 64'd90291986432, - 64'd326352864, 64'd93595976, 64'd2567953973248, - 64'd92239462400, - 64'd215365024, 64'd93990832, 64'd2521365741568, - 64'd94098808832, - 64'd102901504, 64'd94183904, 64'd2473870229504, - 64'd95868690432, 64'd10874321, 64'd94175632, 64'd2425512263680, - 64'd97547862016, 64'd125798456, 64'd93966792, 64'd2376337719296, - 64'd99135217664, 64'd241706592, 64'd93558536, 64'd2326392471552, - 64'd100629733376, 64'd358434368, 64'd92952320, 64'd2275723444224, - 64'd102030532608, 64'd475817568, 64'd92149960, 64'd2224377823232, - 64'd103336837120, 64'd593692416, 64'd91153584, 64'd2172402532352, - 64'd104547975168, 64'd711895808, 64'd89965616, 64'd2119845675008, - 64'd105663406080, 64'd830265472, 64'd88588808, 64'd2066755092480, - 64'd106682703872, 64'd948640384, 64'd87026168, 64'd2013179019264, - 64'd107605540864, 64'd1066860608, 64'd85281016, 64'd1959165689856, - 64'd108431712256, 64'd1184768000, 64'd83356920, 64'd1904763469824, - 64'd109161119744, 64'd1302206208, 64'd81257720, 64'd1850020724736, - 64'd109793796096, 64'd1419020544, 64'd78987496, 64'd1794985820160, - 64'd110329856000, 64'd1535058816, 64'd76550560, 64'd1739706990592, - 64'd110769553408, 64'd1650171136, 64'd73951456, 64'd1684232208384, - 64'd111113216000, 64'd1764210048, 64'd71194960, 64'd1628609576960, - 64'd111361302528, 64'd1877030784, 64'd68286016, 64'd1572886806528, - 64'd111514378240, 64'd1988491648, 64'd65229784, 64'd1517110951936, - 64'd111573098496, 64'd2098454016, 64'd62031604, 64'd1461329330176, - 64'd111538233344, 64'd2206782464, 64'd58696980, 64'd1405588209664, - 64'd111410634752, 64'd2313344512, 64'd55231580, 64'd1349933989888, - 64'd111191261184, 64'd2418012160, 64'd51641208, 64'd1294412021760, - 64'd110881177600, 64'd2520659968, 64'd47931816, 64'd1239067656192, - 64'd110481530880, 64'd2621167360, 64'd44109480, 64'd1183945195520, - 64'd109993558016, 64'd2719416576, 64'd40180376, 64'd1129088679936, - 64'd109418586112, 64'd2815294720, 64'd36150796, 64'd1074540904448, - 64'd108758032384, 64'd2908692992, 64'd32027118, 64'd1020344598528, - 64'd108013395968, 64'd2999506176, 64'd27815800, 64'd966541312000, - 64'd107186249728, 64'd3087634176, 64'd23523372, 64'd913171808256, - 64'd106278248448, 64'd3172980992, 64'd19156418, 64'd860276260864, - 64'd105291128832, 64'd3255454720, 64'd14721570, 64'd807893598208, - 64'd104226684928, 64'd3334968832, 64'd10225500, 64'd756062093312, - 64'd103086809088, 64'd3411440896, 64'd5674904, 64'd704819036160, - 64'd101873418240, 64'd3484793344, 64'd1076496, 64'd654200602624, - 64'd100588527616, 64'd3554953472, - 64'd3563006, 64'd604242116608, - 64'd99234201600, 64'd3621852928, - 64'd8236886, 64'd554977656832, - 64'd97812545536, 64'd3685428480, - 64'd12938444, 64'd506440384512, - 64'd96325754880, 64'd3745622272, - 64'd17661002, 64'd458662379520, - 64'd94776033280, 64'd3802380288, - 64'd22397912, 64'd411674476544, - 64'd93165666304, 64'd3855654400, - 64'd27142574, 64'd365506428928, - 64'd91496964096, 64'd3905400576, - 64'd31888434, 64'd320186843136, - 64'd89772285952, 64'd3951580160, - 64'd36628996, 64'd275743080448, - 64'd87994023936, 64'd3994159360, - 64'd41357844, 64'd232201338880, - 64'd86164611072, 64'd4033108992, - 64'd46068624, 64'd189586587648, - 64'd84286504960, 64'd4068405248, - 64'd50755072, 64'd147922534400, - 64'd82362204160, 64'd4100028672, - 64'd55411020, 64'd107231666176, - 64'd80394207232, 64'd4127964928, - 64'd60030396, 64'd67535187968, - 64'd78385053696, 64'd4152204288, - 64'd64607236, 64'd28853045248, - 64'd76337299456, 64'd4172742144, - 64'd69135696, - 64'd8796102656, - 64'd74253508608, 64'd4189577728, - 64'd73610040, - 64'd45394882560, - 64'd72136261632, 64'd4202715904, - 64'd78024672, - 64'd80927219712, - 64'd69988139008, 64'd4212165376, - 64'd82374128, - 64'd115378307072, - 64'd67811745792, 64'd4217939712, - 64'd86653072, - 64'd148734672896, - 64'd65609662464, 64'd4220057088, - 64'd90856336, - 64'd180984119296, - 64'd63384489984, 64'd4218539520, - 64'd94978888, - 64'd212115750912, - 64'd61138817024, 64'd4213413888, - 64'd99015848, - 64'd242119950336, - 64'd58875224064, 64'd4204710912, - 64'd102962496, - 64'd270988410880, - 64'd56596283392, 64'd4192465408, - 64'd106814296, - 64'd298714103808, - 64'd54304550912, 64'd4176716800, - 64'd110566872, - 64'd325291245568, - 64'd52002574336, 64'd4157507328, - 64'd114216008, - 64'd350715379712, - 64'd49692868608, 64'd4134884352, - 64'd117757672, - 64'd374983262208, - 64'd47377944576, 64'd4108897792, - 64'd121188032, - 64'd398092861440, - 64'd45060276224, 64'd4079602432, - 64'd124503416, - 64'd420043489280, - 64'd42742312960, 64'd4047055104, - 64'd127700336, - 64'd440835538944, - 64'd40426479616, 64'd4011317248, - 64'd130775512, - 64'd460470714368, - 64'd38115160064, 64'd3972453120, - 64'd133725848, - 64'd478951833600, - 64'd35810713600, 64'd3930530048, - 64'd136548432, - 64'd496282959872, - 64'd33515456512, 64'd3885618688, - 64'd139240544, - 64'd512469204992, - 64'd31231666176, 64'd3837792256, - 64'd141799680, - 64'd527516893184, - 64'd28961583104, 64'd3787126784, - 64'd144223504, - 64'd541433430016, - 64'd26707396608, 64'd3733701376, - 64'd146509920, - 64'd554227335168, - 64'd24471257088, 64'd3677597184, - 64'd148656976, - 64'd565908078592, - 64'd22255263744, 64'd3618898176, - 64'd150662944, - 64'd576486244352, - 64'd20061468672, 64'd3557690112, - 64'd152526320, - 64'd585973563392, - 64'd17891870720, 64'd3494061312, - 64'd154245744, - 64'd594382487552, - 64'd15748417536, 64'd3428102144, - 64'd155820096, - 64'd601726648320, - 64'd13632999424, 64'd3359904000, - 64'd157248432, - 64'd608020463616, - 64'd11547452416, 64'd3289561088, - 64'd158530016, - 64'd613279399936, - 64'd9493555200, 64'd3217168384, - 64'd159664272, - 64'd617519579136, - 64'd7473025536, 64'd3142822912, - 64'd160650880, - 64'd620758237184, - 64'd5487523328, 64'd3066622720, - 64'd161489648, - 64'd623013199872, - 64'd3538644224, 64'd2988666624, - 64'd162180592, - 64'd624303276032, - 64'd1627923072, 64'd2909055232, - 64'd162723920, - 64'd624647733248, 64'd243169680, 64'd2827889664, - 64'd163120048, - 64'd624066887680, 64'd2073228160, 64'd2745271552, - 64'd163369504, - 64'd622581579776, 64'd3860911872, 64'd2661303808, - 64'd163473072, - 64'd620213305344, 64'd5604946432, 64'd2576089088, - 64'd163431664, - 64'd616984084480, 64'd7304124928, 64'd2489731072, - 64'd163246368, - 64'd612916789248, 64'd8957306880, 64'd2402333184, - 64'd162918464, - 64'd608034619392, 64'd10563420160, 64'd2313999360, - 64'd162449360, - 64'd602361430016, 64'd12121461760, 64'd2224832768, - 64'd161840640, - 64'd595921338368, 64'd13630494720, 64'd2134937088, - 64'd161094080, - 64'd588739248128, 64'd15089655808, 64'd2044415744, - 64'd160211552, - 64'd580840128512, 64'd16498144256, 64'd1953371392, - 64'd159195120, - 64'd572249669632, 64'd17855234048, 64'd1861906176, - 64'd158046960, - 64'd562993561600, 64'd19160264704, 64'd1770121856, - 64'd156769424, - 64'd553098149888, 64'd20412645376, 64'd1678119168, - 64'd155364944, - 64'd542589812736, 64'd21611853824, 64'd1585998080, - 64'd153836160, - 64'd531495256064, 64'd22757437440, 64'd1493857408, - 64'd152185744, - 64'd519841382400, 64'd23849011200, 64'd1401795200, - 64'd150416576, - 64'd507655290880, 64'd24886253568, 64'd1309908096, - 64'd148531600, - 64'd494964211712, 64'd25868914688, 64'd1218291200, - 64'd146533888, - 64'd481795506176, 64'd26796810240, 64'd1127038592, - 64'd144426608, - 64'd468176568320, 64'd27669821440, 64'd1036242496, - 64'd142213024, - 64'd454134824960, 64'd28487892992, 64'd945993792, - 64'd139896528, - 64'd439697801216, 64'd29251037184, 64'd856381504, - 64'd137480544, - 64'd424892956672, 64'd29959323648, 64'd767492992, - 64'd134968656, - 64'd409747619840, 64'd30612889600, 64'd679413632, - 64'd132364440, - 64'd394289152000, 64'd31211931648, 64'd592226880, - 64'd129671616, - 64'd378544717824, 64'd31756709888, 64'd506014144, - 64'd126893928, - 64'd362541416448, 64'd32247535616, 64'd420854784, - 64'd124035200, - 64'd346306117632, 64'd32684787712, 64'd336825984, - 64'd121099320, - 64'd329865494528, 64'd33068896256, 64'd254002592, - 64'd118090200, - 64'd313245990912, 64'd33400346624, 64'd172457248, - 64'd115011824, - 64'd296473821184, 64'd33679681536, 64'd92260200, - 64'd111868200, - 64'd279574904832, 64'd33907492864, 64'd13479277, - 64'd108663376, - 64'd262574817280, 64'd34084423680, - 64'd63820176, - 64'd105401440, - 64'd245498839040, 64'd34211174400, - 64'd139575328, - 64'd102086472, - 64'd228371890176, 64'd34288482304, - 64'd213725904, - 64'd98722608, - 64'd211218464768, 64'd34317139968, - 64'd286214240, - 64'd95313960, - 64'd194062712832, 64'd34297980928, - 64'd356985312, - 64'd91864688, - 64'd176928309248, 64'd34231885824, - 64'd425986784, - 64'd88378912, - 64'd159838502912, 64'd34119774208, - 64'd493169024, - 64'd84860784, - 64'd142816051200, 64'd33962604544, - 64'd558485120, - 64'd81314424, - 64'd125883236352, 64'd33761378304, - 64'd621890880, - 64'd77743960, - 64'd109061840896, 64'd33517131776, - 64'd683344960, - 64'd74153472, - 64'd92373098496, 64'd33230934016, - 64'd742808768, - 64'd70547056, - 64'd75837718528, 64'd32903890944, - 64'd800246464, - 64'd66928744, - 64'd59475828736, 64'd32537139200, - 64'd855625088, - 64'd63302560, - 64'd43306999808, 64'd32131840000, - 64'd908914368, - 64'd59672484, - 64'd27350212608, 64'd31689191424, - 64'd960087104, - 64'd56042448, - 64'd11623832576, 64'd31210409984, - 64'd1009118528, - 64'd52416348, 64'd3854381568, 64'd30696738816, - 64'd1055987008, - 64'd48798032, 64'd19067301888, 64'd30149447680, - 64'd1100673536, - 64'd45191280, 64'd33998438400, 64'd29569818624, - 64'd1143161856, - 64'd41599828, 64'd48631947264, 64'd28959158272, - 64'd1183438592, - 64'd38027344, 64'd62952644608, 64'd28318789632, - 64'd1221492864, - 64'd34477432, 64'd76946006016, 64'd27650050048, - 64'd1257316992, - 64'd30953630, 64'd90598187008, 64'd26954289152, - 64'd1290905472, - 64'd27459396, 64'd103896023040, 64'd26232868864, - 64'd1322255616, - 64'd23998120, 64'd116827013120, 64'd25487161344, - 64'd1351367680, - 64'd20573110, 64'd129379360768, 64'd24718544896, - 64'd1378243968, - 64'd17187588, 64'd141541965824, 64'd23928403968, - 64'd1402889856, - 64'd13844698, 64'd153304416256, 64'd23118131200, - 64'd1425313024, - 64'd10547491, 64'd164656971776, 64'd22289115136, - 64'd1445523584, - 64'd7298930, 64'd175590637568, 64'd21442752512, - 64'd1463533952, - 64'd4101886, 64'd186097074176, 64'd20580433920, - 64'd1479359360, - 64'd959131, 64'd196168646656, 64'd19703549952, - 64'd1493017088, 64'd2126656, 64'd205798424576, 64'd18813483008, - 64'd1504526720, 64'd5152898, 64'd214980149248, 64'd17911617536, - 64'd1513909888, 64'd8117120, 64'd223708299264, 64'd16999323648, - 64'd1521190912, 64'd11016947, 64'd231977975808, 64'd16077966336, - 64'd1526395776, 64'd13850111, 64'd239784984576, 64'd15148897280, - 64'd1529552640, 64'd16614449, 64'd247125803008, 64'd14213457920, - 64'd1530691712, 64'd19307906, 64'd253997596672, 64'd13272977408, - 64'd1529845120, 64'd21928534, 64'd260398153728, 64'd12328769536, - 64'd1527046912, 64'd24474498, 64'd266325950464, 64'd11382128640, - 64'd1522332672, 64'd26944068, 64'd271780102144, 64'd10434337792, - 64'd1515740160, 64'd29335628, 64'd276760297472, 64'd9486654464, - 64'd1507308416, 64'd31647676, 64'd281266978816, 64'd8540322304, - 64'd1497078272, 64'd33878816, 64'd285301080064, 64'd7596559872, - 64'd1485092096, 64'd36027768, 64'd288864174080, 64'd6656563712, - 64'd1471393536, 64'd38093364, 64'd291958456320, 64'd5721507840, - 64'd1456027776, 64'd40074548, 64'd294586679296, 64'd4792541184, - 64'd1439041408, 64'd41970372, 64'd296752185344, 64'd3870787072, - 64'd1420482048, 64'd43780008, 64'd298458841088, 64'd2957342208, - 64'd1400398592, 64'd45502732, 64'd299711102976, 64'd2053275520, - 64'd1378840960, 64'd47137936, 64'd300513853440, 64'd1159627392, - 64'd1355860096, 64'd48685116, 64'd300872630272, 64'd277409216, - 64'd1331507840, 64'd50143884, 64'd300793331712, - 64'd592398208, - 64'd1305837056, 64'd51513952, 64'd300282445824, - 64'd1448844928, - 64'd1278901376, 64'd52795148, 64'd299346886656, - 64'd2291012352, - 64'd1250754816, 64'd53987404, 64'd297993961472, - 64'd3118014208, - 64'd1221452416, 64'd55090748, 64'd296231534592, - 64'd3928997632, - 64'd1191049728, 64'd56105320, 64'd294067798016, - 64'd4723142656, - 64'd1159602560, 64'd57031364, 64'd291511336960, - 64'd5499663360, - 64'd1127167232, 64'd57869220, 64'd288571195392, - 64'd6257808896, - 64'd1093800576, 64'd58619320, 64'd285256712192, - 64'd6996861440, - 64'd1059559552, 64'd59282200, 64'd281577619456, - 64'd7716141056, - 64'd1024501184, 64'd59858492, 64'd277543976960, - 64'd8415001088, - 64'd988682816, 64'd60348920, 64'd273166123008, - 64'd9092832256, - 64'd952161856, 64'd60754288, 64'd268454739968, - 64'd9749059584, - 64'd914995456, 64'd61075508, 64'd263420755968, - 64'd10383145984, - 64'd877240960, 64'd61313560, 64'd258075361280, - 64'd10994589696, - 64'd838955392, 64'd61469516, 64'd252430008320, - 64'd11582924800, - 64'd800195648, 64'd61544524, 64'd246496362496, - 64'd12147724288, - 64'd761018176, 64'd61539824, 64'd240286269440, - 64'd12688594944, - 64'd721479296, 64'd61456716, 64'd233811820544, - 64'd13205181440, - 64'd681634752, 64'd61296580, 64'd227085189120, - 64'd13697163264, - 64'd641539776, 64'd61060876, 64'd220118794240, - 64'd14164257792, - 64'd601249280, 64'd60751116, 64'd212925120512, - 64'd14606216192, - 64'd560817408, 64'd60368888, 64'd205516800000, - 64'd15022828544, - 64'd520297600, 64'd59915840, 64'd197906546688, - 64'd15413916672, - 64'd479742752, 64'd59393688, 64'd190107172864, - 64'd15779340288, - 64'd439204928, 64'd58804188, 64'd182131507200, - 64'd16118992896, - 64'd398735328, 64'd58149164, 64'd173992476672, - 64'd16432802816, - 64'd358384352, 64'd57430484, 64'd165703024640, - 64'd16720731136, - 64'd318201440, 64'd56650076, 64'd157276061696, - 64'd16982773760, - 64'd278235136, 64'd55809896, 64'd148724563968, - 64'd17218959360, - 64'd238532896, 64'd54911956, 64'd140061409280, - 64'd17429350400, - 64'd199141184, 64'd53958296, 64'd131299491840, - 64'd17614036992, - 64'd160105344, 64'd52951008, 64'd122451632128, - 64'd17773146112, - 64'd121469616, 64'd51892204, 64'd113530585088, - 64'd17906831360, - 64'd83277048, 64'd50784028, 64'd104549007360, - 64'd18015279104, - 64'd45569488, 64'd49628656, 64'd95519473664, - 64'd18098704384, - 64'd8387556, 64'd48428288, 64'd86454435840, - 64'd18157350912, 64'd28229402, 64'd47185140, 64'd77366206464, - 64'd18191486976, 64'd64243336, 64'd45901452, 64'd68266983424, - 64'd18201415680, 64'd99617528, 64'd44579476, 64'd59168776192, - 64'd18187460608, 64'd134316608, 64'd43221476, 64'd50083442688, - 64'd18149971968, 64'd168306576, 64'd41829732, 64'd41022660608, - 64'd18089326592, 64'd201554848, 64'd40406520, 64'd31997908992, - 64'd18005925888, 64'd234030224, 64'd38954128, 64'd23020460032, - 64'd17900189696, 64'd265702976, 64'd37474844, 64'd14101369856, - 64'd17772564480, 64'd296544800, 64'd35970948, 64'd5251466752, - 64'd17623517184, 64'd326528896, 64'd34444728, - 64'd3518658560, - 64'd17453537280, 64'd355629856, 64'd32898450, - 64'd12198665216, - 64'd17263128576, 64'd383823840, 64'd31334380, - 64'd20778469376, - 64'd17052819456, 64'd411088448, 64'd29754768, - 64'd29248258048, - 64'd16823151616, 64'd437402848, 64'd28161850, - 64'd37598486528, - 64'd16574686208, 64'd462747616, 64'd26557844, - 64'd45819908096, - 64'd16307999744, 64'd487104896, 64'd24944950, - 64'd53903548416, - 64'd16023682048, 64'd510458336, 64'd23325340, - 64'd61840748544, - 64'd15722339328, 64'd532793056, 64'd21701168, - 64'd69623152640, - 64'd15404589056, 64'd554095680, 64'd20074556, - 64'd77242712064, - 64'd15071063040, 64'd574354368, 64'd18447600, - 64'd84691689472, - 64'd14722400256, 64'd593558656, 64'd16822366, - 64'd91962695680, - 64'd14359252992, 64'd611699712, 64'd15200882, - 64'd99048644608, - 64'd13982282752, 64'd628770112, 64'd13585143, - 64'd105942786048, - 64'd13592156160, 64'd644763840, 64'd11977109, - 64'd112638713856, - 64'd13189551104, 64'd659676288, 64'd10378697, - 64'd119130365952, - 64'd12775148544, 64'd673504448, 64'd8791785, - 64'd125412016128, - 64'd12349637632, 64'd686246528, 64'd7218210, - 64'd131478265856, - 64'd11913708544, 64'd697902208, 64'd5659761, - 64'd137324101632, - 64'd11468056576, 64'd708472576, 64'd4118186, - 64'd142944829440, - 64'd11013382144, 64'd717960064, 64'd2595181, - 64'd148336099328, - 64'd10550381568, 64'd726368320, 64'd1092397, - 64'd153493929984, - 64'd10079757312, 64'd733702400, - 64'd388567, - 64'd158414700544, - 64'd9602208768, 64'd739968640, - 64'd1846161, - 64'd163095101440, - 64'd9118435328, 64'd745174528, - 64'd3278891, - 64'd167532216320, - 64'd8629133312, 64'd749328960, - 64'd4685312, - 64'd171723423744, - 64'd8134998016, 64'd752441856, - 64'd6064036, - 64'd175666511872, - 64'd7636720128, 64'd754524288, - 64'd7413731, - 64'd179359580160, - 64'd7134985728, 64'd755588608, - 64'd8733119, - 64'd182801039360, - 64'd6630476288, 64'd755648192, - 64'd10020980, - 64'd185989693440, - 64'd6123866624, 64'd754717504, - 64'd11276151, - 64'd188924674048, - 64'd5615825408, 64'd752811968, - 64'd12497527, - 64'd191605391360, - 64'd5107013632, 64'd749948096, - 64'd13684064, - 64'd194031665152, - 64'd4598084096, 64'd746143296, - 64'd14834774, - 64'd196203560960, - 64'd4089680640, 64'd741416064, - 64'd15948730, - 64'd198121537536, - 64'd3582437376, 64'd735785600, - 64'd17025066, - 64'd199786299392, - 64'd3076978176, 64'd729272064, - 64'd18062970, - 64'd201198911488, - 64'd2573916416, 64'd721896384, - 64'd19061700, - 64'd202360717312, - 64'd2073853440, 64'd713680384, - 64'd20020564, - 64'd203273371648, - 64'd1577378816, 64'd704646400, - 64'd20938938, - 64'd203938791424, - 64'd1085069056, 64'd694817792, - 64'd21816254, - 64'd204359221248, - 64'd597488000, 64'd684218240, - 64'd22652002, - 64'd204537151488, - 64'd115185360, 64'd672872384, - 64'd23445736, - 64'd204475383808, 64'd361303328, 64'd660805248, - 64'd24197068, - 64'd204176916480, 64'd831457152, 64'd648042368, - 64'd24905666, - 64'd203645059072, 64'd1294770432, 64'd634609984, - 64'd25571260, - 64'd202883366912, 64'd1750752896, 64'd620534592, - 64'd26193636, - 64'd201895608320, 64'd2198930432, 64'd605843264, - 64'd26772638, - 64'd200685813760, 64'd2638845440, 64'd590563392, - 64'd27308166, - 64'd199258210304, 64'd3070056448, 64'd574722752, - 64'd27800178, - 64'd197617270784, 64'd3492139264, 64'd558349440, - 64'd28248684, - 64'd195767664640, 64'd3904687104, 64'd541471680, - 64'd28653752, - 64'd193714241536, 64'd4307311104, 64'd524118112, - 64'd29015500};

	localparam logic signed[63:0] hb[0:1199] = {64'd3360891076608, 64'd1740072192, - 64'd2258560256, - 64'd2309433, 64'd3359151226880, 64'd5218416128, - 64'd2253798656, - 64'd6921711, 64'd3355673624576, 64'd8691364864, - 64'd2244285696, - 64'd11514461, 64'd3350461415424, 64'd12155332608, - 64'd2230039808, - 64'd16075163, 64'd3343520366592, 64'd15606747136, - 64'd2211088640, - 64'd20591730, 64'd3334857293824, 64'd19042058240, - 64'd2187467776, - 64'd25052516, 64'd3324481372160, 64'd22457741312, - 64'd2159221248, - 64'd29446316, 64'd3312403349504, 64'd25850302464, - 64'd2126401536, - 64'd33762368, 64'd3298635546624, 64'd29216280576, - 64'd2089067776, - 64'd37990368, 64'd3283192119296, 64'd32552259584, - 64'd2047287168, - 64'd42120460, 64'd3266088796160, 64'd35854868480, - 64'd2001134208, - 64'd46143240, 64'd3247343403008, 64'd39120789504, - 64'd1950690048, - 64'd50049756, 64'd3226974814208, 64'd42346749952, - 64'd1896042368, - 64'd53831528, 64'd3205003739136, 64'd45529546752, - 64'd1837285632, - 64'd57480512, 64'd3181452984320, 64'd48666038272, - 64'd1774520192, - 64'd60989140, 64'd3156345880576, 64'd51753148416, - 64'd1707852160, - 64'd64350292, 64'd3129708380160, 64'd54787874816, - 64'd1637393280, - 64'd67557296, 64'd3101567221760, 64'd57767292928, - 64'd1563260672, - 64'd70603936, 64'd3071950979072, 64'd60688547840, - 64'd1485576448, - 64'd73484464, 64'd3040889012224, 64'd63548878848, - 64'd1404467200, - 64'd76193552, 64'd3008412516352, 64'd66345603072, - 64'd1320064256, - 64'd78726344, 64'd2974554259456, 64'd69076131840, - 64'd1232503040, - 64'd81078400, 64'd2939347795968, 64'd71737966592, - 64'd1141922688, - 64'd83245736, 64'd2902828253184, 64'd74328702976, - 64'd1048465984, - 64'd85224800, 64'd2865031544832, 64'd76846030848, - 64'd952279104, - 64'd87012456, 64'd2825994895360, 64'd79287738368, - 64'd853511232, - 64'd88605992, 64'd2785756577792, 64'd81651720192, - 64'd752314240, - 64'd90003120, 64'd2744356438016, 64'd83935985664, - 64'd648842368, - 64'd91201968, 64'd2701834321920, 64'd86138626048, - 64'd543252352, - 64'd92201048, 64'd2658231648256, 64'd88257855488, - 64'd435702464, - 64'd92999280, 64'd2613590622208, 64'd90291986432, - 64'd326352864, - 64'd93595976, 64'd2567953973248, 64'd92239462400, - 64'd215365024, - 64'd93990832, 64'd2521365741568, 64'd94098808832, - 64'd102901504, - 64'd94183904, 64'd2473870229504, 64'd95868690432, 64'd10874321, - 64'd94175632, 64'd2425512263680, 64'd97547862016, 64'd125798456, - 64'd93966792, 64'd2376337719296, 64'd99135217664, 64'd241706592, - 64'd93558536, 64'd2326392471552, 64'd100629733376, 64'd358434368, - 64'd92952320, 64'd2275723444224, 64'd102030532608, 64'd475817568, - 64'd92149960, 64'd2224377823232, 64'd103336837120, 64'd593692416, - 64'd91153584, 64'd2172402532352, 64'd104547975168, 64'd711895808, - 64'd89965616, 64'd2119845675008, 64'd105663406080, 64'd830265472, - 64'd88588808, 64'd2066755092480, 64'd106682703872, 64'd948640384, - 64'd87026168, 64'd2013179019264, 64'd107605540864, 64'd1066860608, - 64'd85281016, 64'd1959165689856, 64'd108431712256, 64'd1184768000, - 64'd83356920, 64'd1904763469824, 64'd109161119744, 64'd1302206208, - 64'd81257720, 64'd1850020724736, 64'd109793796096, 64'd1419020544, - 64'd78987496, 64'd1794985820160, 64'd110329856000, 64'd1535058816, - 64'd76550560, 64'd1739706990592, 64'd110769553408, 64'd1650171136, - 64'd73951456, 64'd1684232208384, 64'd111113216000, 64'd1764210048, - 64'd71194960, 64'd1628609576960, 64'd111361302528, 64'd1877030784, - 64'd68286016, 64'd1572886806528, 64'd111514378240, 64'd1988491648, - 64'd65229784, 64'd1517110951936, 64'd111573098496, 64'd2098454016, - 64'd62031604, 64'd1461329330176, 64'd111538233344, 64'd2206782464, - 64'd58696980, 64'd1405588209664, 64'd111410634752, 64'd2313344512, - 64'd55231580, 64'd1349933989888, 64'd111191261184, 64'd2418012160, - 64'd51641208, 64'd1294412021760, 64'd110881177600, 64'd2520659968, - 64'd47931816, 64'd1239067656192, 64'd110481530880, 64'd2621167360, - 64'd44109480, 64'd1183945195520, 64'd109993558016, 64'd2719416576, - 64'd40180376, 64'd1129088679936, 64'd109418586112, 64'd2815294720, - 64'd36150796, 64'd1074540904448, 64'd108758032384, 64'd2908692992, - 64'd32027118, 64'd1020344598528, 64'd108013395968, 64'd2999506176, - 64'd27815800, 64'd966541312000, 64'd107186249728, 64'd3087634176, - 64'd23523372, 64'd913171808256, 64'd106278248448, 64'd3172980992, - 64'd19156418, 64'd860276260864, 64'd105291128832, 64'd3255454720, - 64'd14721570, 64'd807893598208, 64'd104226684928, 64'd3334968832, - 64'd10225500, 64'd756062093312, 64'd103086809088, 64'd3411440896, - 64'd5674904, 64'd704819036160, 64'd101873418240, 64'd3484793344, - 64'd1076496, 64'd654200602624, 64'd100588527616, 64'd3554953472, 64'd3563006, 64'd604242116608, 64'd99234201600, 64'd3621852928, 64'd8236886, 64'd554977656832, 64'd97812545536, 64'd3685428480, 64'd12938444, 64'd506440384512, 64'd96325754880, 64'd3745622272, 64'd17661002, 64'd458662379520, 64'd94776033280, 64'd3802380288, 64'd22397912, 64'd411674476544, 64'd93165666304, 64'd3855654400, 64'd27142574, 64'd365506428928, 64'd91496964096, 64'd3905400576, 64'd31888434, 64'd320186843136, 64'd89772285952, 64'd3951580160, 64'd36628996, 64'd275743080448, 64'd87994023936, 64'd3994159360, 64'd41357844, 64'd232201338880, 64'd86164611072, 64'd4033108992, 64'd46068624, 64'd189586587648, 64'd84286504960, 64'd4068405248, 64'd50755072, 64'd147922534400, 64'd82362204160, 64'd4100028672, 64'd55411020, 64'd107231666176, 64'd80394207232, 64'd4127964928, 64'd60030396, 64'd67535187968, 64'd78385053696, 64'd4152204288, 64'd64607236, 64'd28853045248, 64'd76337299456, 64'd4172742144, 64'd69135696, - 64'd8796102656, 64'd74253508608, 64'd4189577728, 64'd73610040, - 64'd45394882560, 64'd72136261632, 64'd4202715904, 64'd78024672, - 64'd80927219712, 64'd69988139008, 64'd4212165376, 64'd82374128, - 64'd115378307072, 64'd67811745792, 64'd4217939712, 64'd86653072, - 64'd148734672896, 64'd65609662464, 64'd4220057088, 64'd90856336, - 64'd180984119296, 64'd63384489984, 64'd4218539520, 64'd94978888, - 64'd212115750912, 64'd61138817024, 64'd4213413888, 64'd99015848, - 64'd242119950336, 64'd58875224064, 64'd4204710912, 64'd102962496, - 64'd270988410880, 64'd56596283392, 64'd4192465408, 64'd106814296, - 64'd298714103808, 64'd54304550912, 64'd4176716800, 64'd110566872, - 64'd325291245568, 64'd52002574336, 64'd4157507328, 64'd114216008, - 64'd350715379712, 64'd49692868608, 64'd4134884352, 64'd117757672, - 64'd374983262208, 64'd47377944576, 64'd4108897792, 64'd121188032, - 64'd398092861440, 64'd45060276224, 64'd4079602432, 64'd124503416, - 64'd420043489280, 64'd42742312960, 64'd4047055104, 64'd127700336, - 64'd440835538944, 64'd40426479616, 64'd4011317248, 64'd130775512, - 64'd460470714368, 64'd38115160064, 64'd3972453120, 64'd133725848, - 64'd478951833600, 64'd35810713600, 64'd3930530048, 64'd136548432, - 64'd496282959872, 64'd33515456512, 64'd3885618688, 64'd139240544, - 64'd512469204992, 64'd31231666176, 64'd3837792256, 64'd141799680, - 64'd527516893184, 64'd28961583104, 64'd3787126784, 64'd144223504, - 64'd541433430016, 64'd26707396608, 64'd3733701376, 64'd146509920, - 64'd554227335168, 64'd24471257088, 64'd3677597184, 64'd148656976, - 64'd565908078592, 64'd22255263744, 64'd3618898176, 64'd150662944, - 64'd576486244352, 64'd20061468672, 64'd3557690112, 64'd152526320, - 64'd585973563392, 64'd17891870720, 64'd3494061312, 64'd154245744, - 64'd594382487552, 64'd15748417536, 64'd3428102144, 64'd155820096, - 64'd601726648320, 64'd13632999424, 64'd3359904000, 64'd157248432, - 64'd608020463616, 64'd11547452416, 64'd3289561088, 64'd158530016, - 64'd613279399936, 64'd9493555200, 64'd3217168384, 64'd159664272, - 64'd617519579136, 64'd7473025536, 64'd3142822912, 64'd160650880, - 64'd620758237184, 64'd5487523328, 64'd3066622720, 64'd161489648, - 64'd623013199872, 64'd3538644224, 64'd2988666624, 64'd162180592, - 64'd624303276032, 64'd1627923072, 64'd2909055232, 64'd162723920, - 64'd624647733248, - 64'd243169680, 64'd2827889664, 64'd163120048, - 64'd624066887680, - 64'd2073228160, 64'd2745271552, 64'd163369504, - 64'd622581579776, - 64'd3860911872, 64'd2661303808, 64'd163473072, - 64'd620213305344, - 64'd5604946432, 64'd2576089088, 64'd163431664, - 64'd616984084480, - 64'd7304124928, 64'd2489731072, 64'd163246368, - 64'd612916789248, - 64'd8957306880, 64'd2402333184, 64'd162918464, - 64'd608034619392, - 64'd10563420160, 64'd2313999360, 64'd162449360, - 64'd602361430016, - 64'd12121461760, 64'd2224832768, 64'd161840640, - 64'd595921338368, - 64'd13630494720, 64'd2134937088, 64'd161094080, - 64'd588739248128, - 64'd15089655808, 64'd2044415744, 64'd160211552, - 64'd580840128512, - 64'd16498144256, 64'd1953371392, 64'd159195120, - 64'd572249669632, - 64'd17855234048, 64'd1861906176, 64'd158046960, - 64'd562993561600, - 64'd19160264704, 64'd1770121856, 64'd156769424, - 64'd553098149888, - 64'd20412645376, 64'd1678119168, 64'd155364944, - 64'd542589812736, - 64'd21611853824, 64'd1585998080, 64'd153836160, - 64'd531495256064, - 64'd22757437440, 64'd1493857408, 64'd152185744, - 64'd519841382400, - 64'd23849011200, 64'd1401795200, 64'd150416576, - 64'd507655290880, - 64'd24886253568, 64'd1309908096, 64'd148531600, - 64'd494964211712, - 64'd25868914688, 64'd1218291200, 64'd146533888, - 64'd481795506176, - 64'd26796810240, 64'd1127038592, 64'd144426608, - 64'd468176568320, - 64'd27669821440, 64'd1036242496, 64'd142213024, - 64'd454134824960, - 64'd28487892992, 64'd945993792, 64'd139896528, - 64'd439697801216, - 64'd29251037184, 64'd856381504, 64'd137480544, - 64'd424892956672, - 64'd29959323648, 64'd767492992, 64'd134968656, - 64'd409747619840, - 64'd30612889600, 64'd679413632, 64'd132364440, - 64'd394289152000, - 64'd31211931648, 64'd592226880, 64'd129671616, - 64'd378544717824, - 64'd31756709888, 64'd506014144, 64'd126893928, - 64'd362541416448, - 64'd32247535616, 64'd420854784, 64'd124035200, - 64'd346306117632, - 64'd32684787712, 64'd336825984, 64'd121099320, - 64'd329865494528, - 64'd33068896256, 64'd254002592, 64'd118090200, - 64'd313245990912, - 64'd33400346624, 64'd172457248, 64'd115011824, - 64'd296473821184, - 64'd33679681536, 64'd92260200, 64'd111868200, - 64'd279574904832, - 64'd33907492864, 64'd13479277, 64'd108663376, - 64'd262574817280, - 64'd34084423680, - 64'd63820176, 64'd105401440, - 64'd245498839040, - 64'd34211174400, - 64'd139575328, 64'd102086472, - 64'd228371890176, - 64'd34288482304, - 64'd213725904, 64'd98722608, - 64'd211218464768, - 64'd34317139968, - 64'd286214240, 64'd95313960, - 64'd194062712832, - 64'd34297980928, - 64'd356985312, 64'd91864688, - 64'd176928309248, - 64'd34231885824, - 64'd425986784, 64'd88378912, - 64'd159838502912, - 64'd34119774208, - 64'd493169024, 64'd84860784, - 64'd142816051200, - 64'd33962604544, - 64'd558485120, 64'd81314424, - 64'd125883236352, - 64'd33761378304, - 64'd621890880, 64'd77743960, - 64'd109061840896, - 64'd33517131776, - 64'd683344960, 64'd74153472, - 64'd92373098496, - 64'd33230934016, - 64'd742808768, 64'd70547056, - 64'd75837718528, - 64'd32903890944, - 64'd800246464, 64'd66928744, - 64'd59475828736, - 64'd32537139200, - 64'd855625088, 64'd63302560, - 64'd43306999808, - 64'd32131840000, - 64'd908914368, 64'd59672484, - 64'd27350212608, - 64'd31689191424, - 64'd960087104, 64'd56042448, - 64'd11623832576, - 64'd31210409984, - 64'd1009118528, 64'd52416348, 64'd3854381568, - 64'd30696738816, - 64'd1055987008, 64'd48798032, 64'd19067301888, - 64'd30149447680, - 64'd1100673536, 64'd45191280, 64'd33998438400, - 64'd29569818624, - 64'd1143161856, 64'd41599828, 64'd48631947264, - 64'd28959158272, - 64'd1183438592, 64'd38027344, 64'd62952644608, - 64'd28318789632, - 64'd1221492864, 64'd34477432, 64'd76946006016, - 64'd27650050048, - 64'd1257316992, 64'd30953630, 64'd90598187008, - 64'd26954289152, - 64'd1290905472, 64'd27459396, 64'd103896023040, - 64'd26232868864, - 64'd1322255616, 64'd23998120, 64'd116827013120, - 64'd25487161344, - 64'd1351367680, 64'd20573110, 64'd129379360768, - 64'd24718544896, - 64'd1378243968, 64'd17187588, 64'd141541965824, - 64'd23928403968, - 64'd1402889856, 64'd13844698, 64'd153304416256, - 64'd23118131200, - 64'd1425313024, 64'd10547491, 64'd164656971776, - 64'd22289115136, - 64'd1445523584, 64'd7298930, 64'd175590637568, - 64'd21442752512, - 64'd1463533952, 64'd4101886, 64'd186097074176, - 64'd20580433920, - 64'd1479359360, 64'd959131, 64'd196168646656, - 64'd19703549952, - 64'd1493017088, - 64'd2126656, 64'd205798424576, - 64'd18813483008, - 64'd1504526720, - 64'd5152898, 64'd214980149248, - 64'd17911617536, - 64'd1513909888, - 64'd8117120, 64'd223708299264, - 64'd16999323648, - 64'd1521190912, - 64'd11016947, 64'd231977975808, - 64'd16077966336, - 64'd1526395776, - 64'd13850111, 64'd239784984576, - 64'd15148897280, - 64'd1529552640, - 64'd16614449, 64'd247125803008, - 64'd14213457920, - 64'd1530691712, - 64'd19307906, 64'd253997596672, - 64'd13272977408, - 64'd1529845120, - 64'd21928534, 64'd260398153728, - 64'd12328769536, - 64'd1527046912, - 64'd24474498, 64'd266325950464, - 64'd11382128640, - 64'd1522332672, - 64'd26944068, 64'd271780102144, - 64'd10434337792, - 64'd1515740160, - 64'd29335628, 64'd276760297472, - 64'd9486654464, - 64'd1507308416, - 64'd31647676, 64'd281266978816, - 64'd8540322304, - 64'd1497078272, - 64'd33878816, 64'd285301080064, - 64'd7596559872, - 64'd1485092096, - 64'd36027768, 64'd288864174080, - 64'd6656563712, - 64'd1471393536, - 64'd38093364, 64'd291958456320, - 64'd5721507840, - 64'd1456027776, - 64'd40074548, 64'd294586679296, - 64'd4792541184, - 64'd1439041408, - 64'd41970372, 64'd296752185344, - 64'd3870787072, - 64'd1420482048, - 64'd43780008, 64'd298458841088, - 64'd2957342208, - 64'd1400398592, - 64'd45502732, 64'd299711102976, - 64'd2053275520, - 64'd1378840960, - 64'd47137936, 64'd300513853440, - 64'd1159627392, - 64'd1355860096, - 64'd48685116, 64'd300872630272, - 64'd277409216, - 64'd1331507840, - 64'd50143884, 64'd300793331712, 64'd592398208, - 64'd1305837056, - 64'd51513952, 64'd300282445824, 64'd1448844928, - 64'd1278901376, - 64'd52795148, 64'd299346886656, 64'd2291012352, - 64'd1250754816, - 64'd53987404, 64'd297993961472, 64'd3118014208, - 64'd1221452416, - 64'd55090748, 64'd296231534592, 64'd3928997632, - 64'd1191049728, - 64'd56105320, 64'd294067798016, 64'd4723142656, - 64'd1159602560, - 64'd57031364, 64'd291511336960, 64'd5499663360, - 64'd1127167232, - 64'd57869220, 64'd288571195392, 64'd6257808896, - 64'd1093800576, - 64'd58619320, 64'd285256712192, 64'd6996861440, - 64'd1059559552, - 64'd59282200, 64'd281577619456, 64'd7716141056, - 64'd1024501184, - 64'd59858492, 64'd277543976960, 64'd8415001088, - 64'd988682816, - 64'd60348920, 64'd273166123008, 64'd9092832256, - 64'd952161856, - 64'd60754288, 64'd268454739968, 64'd9749059584, - 64'd914995456, - 64'd61075508, 64'd263420755968, 64'd10383145984, - 64'd877240960, - 64'd61313560, 64'd258075361280, 64'd10994589696, - 64'd838955392, - 64'd61469516, 64'd252430008320, 64'd11582924800, - 64'd800195648, - 64'd61544524, 64'd246496362496, 64'd12147724288, - 64'd761018176, - 64'd61539824, 64'd240286269440, 64'd12688594944, - 64'd721479296, - 64'd61456716, 64'd233811820544, 64'd13205181440, - 64'd681634752, - 64'd61296580, 64'd227085189120, 64'd13697163264, - 64'd641539776, - 64'd61060876, 64'd220118794240, 64'd14164257792, - 64'd601249280, - 64'd60751116, 64'd212925120512, 64'd14606216192, - 64'd560817408, - 64'd60368888, 64'd205516800000, 64'd15022828544, - 64'd520297600, - 64'd59915840, 64'd197906546688, 64'd15413916672, - 64'd479742752, - 64'd59393688, 64'd190107172864, 64'd15779340288, - 64'd439204928, - 64'd58804188, 64'd182131507200, 64'd16118992896, - 64'd398735328, - 64'd58149164, 64'd173992476672, 64'd16432802816, - 64'd358384352, - 64'd57430484, 64'd165703024640, 64'd16720731136, - 64'd318201440, - 64'd56650076, 64'd157276061696, 64'd16982773760, - 64'd278235136, - 64'd55809896, 64'd148724563968, 64'd17218959360, - 64'd238532896, - 64'd54911956, 64'd140061409280, 64'd17429350400, - 64'd199141184, - 64'd53958296, 64'd131299491840, 64'd17614036992, - 64'd160105344, - 64'd52951008, 64'd122451632128, 64'd17773146112, - 64'd121469616, - 64'd51892204, 64'd113530585088, 64'd17906831360, - 64'd83277048, - 64'd50784028, 64'd104549007360, 64'd18015279104, - 64'd45569488, - 64'd49628656, 64'd95519473664, 64'd18098704384, - 64'd8387556, - 64'd48428288, 64'd86454435840, 64'd18157350912, 64'd28229402, - 64'd47185140, 64'd77366206464, 64'd18191486976, 64'd64243336, - 64'd45901452, 64'd68266983424, 64'd18201415680, 64'd99617528, - 64'd44579476, 64'd59168776192, 64'd18187460608, 64'd134316608, - 64'd43221476, 64'd50083442688, 64'd18149971968, 64'd168306576, - 64'd41829732, 64'd41022660608, 64'd18089326592, 64'd201554848, - 64'd40406520, 64'd31997908992, 64'd18005925888, 64'd234030224, - 64'd38954128, 64'd23020460032, 64'd17900189696, 64'd265702976, - 64'd37474844, 64'd14101369856, 64'd17772564480, 64'd296544800, - 64'd35970948, 64'd5251466752, 64'd17623517184, 64'd326528896, - 64'd34444728, - 64'd3518658560, 64'd17453537280, 64'd355629856, - 64'd32898450, - 64'd12198665216, 64'd17263128576, 64'd383823840, - 64'd31334380, - 64'd20778469376, 64'd17052819456, 64'd411088448, - 64'd29754768, - 64'd29248258048, 64'd16823151616, 64'd437402848, - 64'd28161850, - 64'd37598486528, 64'd16574686208, 64'd462747616, - 64'd26557844, - 64'd45819908096, 64'd16307999744, 64'd487104896, - 64'd24944950, - 64'd53903548416, 64'd16023682048, 64'd510458336, - 64'd23325340, - 64'd61840748544, 64'd15722339328, 64'd532793056, - 64'd21701168, - 64'd69623152640, 64'd15404589056, 64'd554095680, - 64'd20074556, - 64'd77242712064, 64'd15071063040, 64'd574354368, - 64'd18447600, - 64'd84691689472, 64'd14722400256, 64'd593558656, - 64'd16822366, - 64'd91962695680, 64'd14359252992, 64'd611699712, - 64'd15200882, - 64'd99048644608, 64'd13982282752, 64'd628770112, - 64'd13585143, - 64'd105942786048, 64'd13592156160, 64'd644763840, - 64'd11977109, - 64'd112638713856, 64'd13189551104, 64'd659676288, - 64'd10378697, - 64'd119130365952, 64'd12775148544, 64'd673504448, - 64'd8791785, - 64'd125412016128, 64'd12349637632, 64'd686246528, - 64'd7218210, - 64'd131478265856, 64'd11913708544, 64'd697902208, - 64'd5659761, - 64'd137324101632, 64'd11468056576, 64'd708472576, - 64'd4118186, - 64'd142944829440, 64'd11013382144, 64'd717960064, - 64'd2595181, - 64'd148336099328, 64'd10550381568, 64'd726368320, - 64'd1092397, - 64'd153493929984, 64'd10079757312, 64'd733702400, 64'd388567, - 64'd158414700544, 64'd9602208768, 64'd739968640, 64'd1846161, - 64'd163095101440, 64'd9118435328, 64'd745174528, 64'd3278891, - 64'd167532216320, 64'd8629133312, 64'd749328960, 64'd4685312, - 64'd171723423744, 64'd8134998016, 64'd752441856, 64'd6064036, - 64'd175666511872, 64'd7636720128, 64'd754524288, 64'd7413731, - 64'd179359580160, 64'd7134985728, 64'd755588608, 64'd8733119, - 64'd182801039360, 64'd6630476288, 64'd755648192, 64'd10020980, - 64'd185989693440, 64'd6123866624, 64'd754717504, 64'd11276151, - 64'd188924674048, 64'd5615825408, 64'd752811968, 64'd12497527, - 64'd191605391360, 64'd5107013632, 64'd749948096, 64'd13684064, - 64'd194031665152, 64'd4598084096, 64'd746143296, 64'd14834774, - 64'd196203560960, 64'd4089680640, 64'd741416064, 64'd15948730, - 64'd198121537536, 64'd3582437376, 64'd735785600, 64'd17025066, - 64'd199786299392, 64'd3076978176, 64'd729272064, 64'd18062970, - 64'd201198911488, 64'd2573916416, 64'd721896384, 64'd19061700, - 64'd202360717312, 64'd2073853440, 64'd713680384, 64'd20020564, - 64'd203273371648, 64'd1577378816, 64'd704646400, 64'd20938938, - 64'd203938791424, 64'd1085069056, 64'd694817792, 64'd21816254, - 64'd204359221248, 64'd597488000, 64'd684218240, 64'd22652002, - 64'd204537151488, 64'd115185360, 64'd672872384, 64'd23445736, - 64'd204475383808, - 64'd361303328, 64'd660805248, 64'd24197068, - 64'd204176916480, - 64'd831457152, 64'd648042368, 64'd24905666, - 64'd203645059072, - 64'd1294770432, 64'd634609984, 64'd25571260, - 64'd202883366912, - 64'd1750752896, 64'd620534592, 64'd26193636, - 64'd201895608320, - 64'd2198930432, 64'd605843264, 64'd26772638, - 64'd200685813760, - 64'd2638845440, 64'd590563392, 64'd27308166, - 64'd199258210304, - 64'd3070056448, 64'd574722752, 64'd27800178, - 64'd197617270784, - 64'd3492139264, 64'd558349440, 64'd28248684, - 64'd195767664640, - 64'd3904687104, 64'd541471680, 64'd28653752, - 64'd193714241536, - 64'd4307311104, 64'd524118112, 64'd29015500};


endpackage
`endif

