// Misc utilities used in several modules

typedef struct packed {
    logic[15:0] r;
    logic[31:16] i;
} complex;