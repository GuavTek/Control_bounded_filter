`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam N = 4;
	localparam COEFF_BIAS = 48;
	localparam logic[63:0] Lfr[0:3] = {277489893271481, 277489893271481, 275315491622285, 275315491622285};
	localparam logic[63:0] Lfi[0:3] = {30020001337947, -30020001337947, 11558098293529, -11558098293529};
	localparam logic[63:0] Lbr[0:3] = {277489893271481, 277489893271481, 275315491622285, 275315491622285};
	localparam logic[63:0] Lbi[0:3] = {30020001337947, -30020001337947, 11558098293529, -11558098293529};
	localparam logic[63:0] Wfr[0:3] = {24193209882, 24193209882, -7887428590, -7887428590};
	localparam logic[63:0] Wfi[0:3] = {29297075841, -29297075841, -33126712469, 33126712469};
	localparam logic[63:0] Wbr[0:3] = {-24193209882, -24193209882, 7887428590, 7887428590};
	localparam logic[63:0] Wbi[0:3] = {-29297075841, 29297075841, 33126712469, -33126712469};
	localparam logic[63:0] Ffr[0:3][0:79] = '{
		'{2678910912348682, 1633669149297615, -134405106412023, -14489081406757, 3471761733289509, 1534935316807140, -154547576200402, -12167341321049, 4211153497515380, 1420087166233641, -172563932222687, -9743629047954, 4889422534499934, 1290723849399400, -188281223922595, -7247706595933, 5499740975037776, 1148585763351890, -201556008143343, -4709673588602, 6036181793402482, 995532040410431, -212275515540637, -2159613203878, 6493772333226378, 833517040657504, -220358442413966, 372755769329, 6868535890318197, 664566135678268, -225755365061278, 2858416831816, 7157521071022570, 490751075721102, -228448778179966, 5269379888993, 7358818790936519, 314165232382821, -228452763163329, 7578988059119, 7471566924126414, 136899005473061, -225812296327788, 9762203913194, 7495942755766966, -38984324020268, -220602211106000, 11795872177577, 7433143529741519, -211472022825834, -212925832011491, 13658956252499, 7285355515665612, -378624356972050, -202913301681643, 15332746247078, 7055712145579892, -538595822537850, -190719625501872, 16801036599608, 6748241887867779, -689654930258371, -176522461172683, 18050271736293, 6367806633571694, -830202339184127, -160519683075600, 19069658617453, 5920031467125635, -958787157130758, -142926753400873, 19851245422781, 5411226778650929, -1074121249927379, -123973933701595, 20389966031699, 4848303747586724, -1175091427164946, -103903371822373, 20683650356549},
		'{2678910912348222, 1633669149297648, -134405106412032, -14489081406755, 3471761733289070, 1534935316807172, -154547576200411, -12167341321048, 4211153497514966, 1420087166233671, -172563932222695, -9743629047952, 4889422534499551, 1290723849399429, -188281223922603, -7247706595932, 5499740975037427, 1148585763351916, -201556008143349, -4709673588600, 6036181793402171, 995532040410455, -212275515540643, -2159613203877, 6493772333226108, 833517040657526, -220358442413972, 372755769330, 6868535890317968, 664566135678286, -225755365061283, 2858416831817, 7157521071022387, 490751075721118, -228448778179969, 5269379888994, 7358818790936382, 314165232382833, -228452763163332, 7578988059119, 7471566924126326, 136899005473070, -225812296327790, 9762203913194, 7495942755766923, -38984324020262, -220602211106001, 11795872177577, 7433143529741523, -211472022825831, -212925832011491, 13658956252499, 7285355515665663, -378624356972050, -202913301681642, 15332746247078, 7055712145579987, -538595822537854, -190719625501870, 16801036599608, 6748241887867917, -689654930258378, -176522461172680, 18050271736292, 6367806633571872, -830202339184137, -160519683075597, 19069658617452, 5920031467125852, -958787157130771, -142926753400869, 19851245422781, 5411226778651180, -1074121249927394, -123973933701590, 20389966031698, 4848303747587006, -1175091427164964, -103903371822367, 20683650356548},
		'{-2621464726625032, -1601298142322358, 114277463862052, -54557765512014, -3402192470904109, -1521613693668172, 101035526953527, -52555428834631, -4143075592769200, -1441949887694716, 88125723066021, -50522608463608, -4844167648167600, -1362478337710847, 75562184921028, -48464973598293, -5505606112696863, -1283363101544773, 63357707642890, -46388011318305, -6127608592847788, -1204760640672868, 51523776702445, -44297022280332, -6710469021379336, -1126819797494854, 40070597533593, -42197116997554, -7254553845722606, -1049681790049648, 29007126689070, -40093212685504, -7760298217955961, -973480223457764, 18341104403946, -37990030657633, -8228202194534652, -898341117369665, 8079088437780, -35892094253348, -8658826953596720, -824382948694780, -1773510931025, -33803727280864, -9052791037303526, -751716708882984, -11212394882364, -31729052956814, -9410766626308762, -680445975029133, -20234339123843, -29671993324251, -9733475853085184, -610666994071677, -28837156170190, -27636269130411, -10021687160474126, -542468779358319, -37019656947170, -25625400145358, -10276211711460314, -475933218855185, -44781611831263, -23642705902492, -10497899855813746, -411135194280852, -52123711232903, -21691306841762, -10687637658882664, -348142710452834, -59047525827614, -19774125836360, -10846343497467206, -287017034141629, -65555466535792, -17893890083631, -10974964727353150, -227812841736200, -71650744348225, -16053133340965},
		'{-2621464726623828, -1601298142322414, 114277463862073, -54557765512018, -3402192470902937, -1521613693668227, 101035526953548, -52555428834635, -4143075592768060, -1441949887694769, 88125723066041, -50522608463611, -4844167648166494, -1362478337710898, 75562184921047, -48464973598296, -5505606112695792, -1283363101544822, 63357707642909, -46388011318308, -6127608592846752, -1204760640672916, 51523776702463, -44297022280336, -6710469021378337, -1126819797494900, 40070597533610, -42197116997558, -7254553845721645, -1049681790049693, 29007126689086, -40093212685508, -7760298217955038, -973480223457806, 18341104403961, -37990030657636, -8228202194533767, -898341117369706, 8079088437795, -35892094253351, -8658826953595873, -824382948694820, -1773510931011, -33803727280867, -9052791037302716, -751716708883021, -11212394882350, -31729052956816, -9410766626307994, -680445975029168, -20234339123830, -29671993324253, -9733475853084454, -610666994071711, -28837156170178, -27636269130413, -10021687160473434, -542468779358351, -37019656947158, -25625400145361, -10276211711459662, -475933218855215, -44781611831252, -23642705902494, -10497899855813134, -411135194280880, -52123711232892, -21691306841764, -10687637658882086, -348142710452861, -59047525827604, -19774125836362, -10846343497466668, -287017034141654, -65555466535783, -17893890083633, -10974964727352650, -227812841736223, -71650744348217, -16053133340967}};
	localparam logic[63:0] Ffi[0:3][0:79] = '{
		'{-7789584925020542, 708887221199158, 206702748225345, -19845819841343, -7393588604643268, 873085743790186, 189441643064671, -21110141804839, -6918639246994867, 1024429359565470, 170276674079435, -22108944360993, -6371556198568730, 1161381434685642, 149461551191332, -22835111110926, -5759879607888508, 1282597644249564, 127264837936302, -23284800600437, -5091771080218742, 1386938313763277, 103966594132111, -23457435961284, -4375908801885497, 1473478185138040, 79854941677750, -23355656937657, -3621378440744956, 1541513537288885, 55222594523002, -22985235482842, -2837561156357778, 1590566623196748, 30363393574268, -22354956512906, -2034020064558232, 1620387416998140, 5568886563156, -21476465781011, -1220386496487038, 1630952695911008, -18875008286193, -20364087183631, -406247372102465, 1622462512239921, -42691217575166, -19034612125145, 398965026813756, 1595334139989243, -65614571842042, -17507063846684, 1186079648425665, 1550193608429831, -87394675671855, -15802439866300, 1946288454422587, 1487864961015521, -107798558746626, -13943435878179, 2671242297735851, 1409357402058381, -126613080816752, -11954154617209, 3353139883456778, 1315850515302490, -143647066875003, -9859803310541, 3984808899006887, 1208677757771555, -158733152334642, -7686383409257, 4559778505553668, 1089308448825112, -171729321708043, -5460376320793, 5072342496187033, 959328488094488, -182520128106280, -3208428846785},
		'{7789584925020678, -708887221199165, -206702748225342, 19845819841342, 7393588604643451, -873085743790196, -189441643064668, 21110141804838, 6918639246995094, -1024429359565484, -170276674079431, 22108944360992, 6371556198568998, -1161381434685658, -149461551191327, 22835111110925, 5759879607888814, -1282597644249583, -127264837936296, 23284800600436, 5091771080219080, -1386938313763298, -103966594132105, 23457435961283, 4375908801885863, -1473478185138064, -79854941677743, 23355656937656, 3621378440745346, -1541513537288910, -55222594522994, 22985235482840, 2837561156358186, -1590566623196775, -30363393574260, 22354956512905, 2034020064558654, -1620387416998168, -5568886563148, 21476465781009, 1220386496487468, -1630952695911038, 18875008286202, 20364087183629, 406247372102900, -1622462512239951, 42691217575174, 19034612125143, -398965026813322, -1595334139989273, 65614571842050, 17507063846682, -1186079648425238, -1550193608429861, 87394675671863, 15802439866299, -1946288454422172, -1487864961015550, 107798558746634, 13943435878177, -2671242297735452, -1409357402058410, 126613080816760, 11954154617207, -3353139883456400, -1315850515302518, 143647066875011, 9859803310540, -3984808899006532, -1208677757771581, 158733152334649, 7686383409256, -4559778505553342, -1089308448825137, 171729321708049, 5460376320792, -5072342496186738, -959328488094511, 182520128106285, 3208428846784},
		'{20410122023596984, -1087203619517777, 261581401330405, -19688353631198, 19855845437227768, -1129165953014674, 260549776479662, -21497800075813, 19281639300793944, -1166937977762846, 258996978016206, -23185429430581, 18689575854732616, -1200612237457261, 256948048973282, -24752655664962, 18081679793730520, -1230286297560720, 254428064696757, -26201094598827, 17459925861202104, -1256062325165291, 251462077212791, -27532552007075, 16826236651983674, -1278046676369314, 248075061960339, -28749011807856, 16182480619338714, -1296349491750649, 244291866905447, -29852624356494, 15530470282089826, -1311084300475151, 240137164048391, -30845694866052, 14871960627433400, -1322367633538259, 235635403329143, -31730671974348, 14208647704754270, -1330318646597064, 230810768931151, -32510136476076, 13542167405539158, -1335058752810478, 225687137978284, -33186790237559, 12874094424288384, -1336711266066034, 220288041614798, -33763445310536, 12205941395145922, -1335401054933668, 214636628453457, -34243013260277, 11539158198806890, -1331254207649389, 208755630372409, -34628494722203, 10875131434119388, -1324397708395326, 202667330637182, -34922969200132, 10215184048673250, -1314959125107046, 196393534320064, -35129585118164, 9560575122561506, -1303066309004502, 189955540985356, -35251550137213, 8912499799410572, -1288847106009427, 183374119605357, -35292121746123, 8272089358702066, -1272429080179444, 176669485668604, -35254598136332},
		'{-20410122023597112, 1087203619517783, -261581401330408, 19688353631199, -19855845437227944, 1129165953014683, -260549776479665, 21497800075814, -19281639300794168, 1166937977762856, -258996978016210, 23185429430582, -18689575854732880, 1200612237457274, -256948048973287, 24752655664963, -18081679793730820, 1230286297560734, -254428064696763, 26201094598828, -17459925861202444, 1256062325165307, -251462077212797, 27532552007076, -16826236651984046, 1278046676369332, -248075061960346, 28749011807857, -16182480619339120, 1296349491750668, -244291866905454, 29852624356495, -15530470282090264, 1311084300475172, -240137164048399, 30845694866053, -14871960627433864, 1322367633538281, -235635403329152, 31730671974350, -14208647704754760, 1330318646597088, -230810768931160, 32510136476078, -13542167405539672, 1335058752810502, -225687137978293, 33186790237561, -12874094424288920, 1336711266066060, -220288041614808, 33763445310538, -12205941395146478, 1335401054933694, -214636628453467, 34243013260279, -11539158198807466, 1331254207649416, -208755630372419, 34628494722205, -10875131434119980, 1324397708395354, -202667330637193, 34922969200134, -10215184048673856, 1314959125107074, -196393534320075, 35129585118166, -9560575122562122, 1303066309004531, -189955540985367, 35251550137215, -8912499799411199, 1288847106009456, -183374119605368, 35292121746125, -8272089358702702, 1272429080179473, -176669485668615, 35254598136334}};
	localparam logic[63:0] Fbr[0:3][0:79] = '{
		'{-2678910912348682, 1633669149297615, 134405106412023, -14489081406757, -3471761733289509, 1534935316807140, 154547576200402, -12167341321049, -4211153497515380, 1420087166233641, 172563932222687, -9743629047954, -4889422534499934, 1290723849399400, 188281223922595, -7247706595933, -5499740975037776, 1148585763351890, 201556008143343, -4709673588602, -6036181793402482, 995532040410431, 212275515540637, -2159613203878, -6493772333226378, 833517040657504, 220358442413966, 372755769329, -6868535890318197, 664566135678268, 225755365061278, 2858416831816, -7157521071022570, 490751075721102, 228448778179966, 5269379888993, -7358818790936519, 314165232382821, 228452763163329, 7578988059119, -7471566924126414, 136899005473061, 225812296327788, 9762203913194, -7495942755766966, -38984324020268, 220602211106000, 11795872177577, -7433143529741519, -211472022825834, 212925832011491, 13658956252499, -7285355515665612, -378624356972050, 202913301681643, 15332746247078, -7055712145579892, -538595822537850, 190719625501872, 16801036599608, -6748241887867779, -689654930258371, 176522461172683, 18050271736293, -6367806633571694, -830202339184127, 160519683075600, 19069658617453, -5920031467125635, -958787157130758, 142926753400873, 19851245422781, -5411226778650929, -1074121249927379, 123973933701595, 20389966031699, -4848303747586724, -1175091427164946, 103903371822373, 20683650356549},
		'{-2678910912348222, 1633669149297648, 134405106412032, -14489081406755, -3471761733289070, 1534935316807172, 154547576200411, -12167341321048, -4211153497514966, 1420087166233671, 172563932222695, -9743629047952, -4889422534499551, 1290723849399429, 188281223922603, -7247706595932, -5499740975037427, 1148585763351916, 201556008143349, -4709673588600, -6036181793402171, 995532040410455, 212275515540643, -2159613203877, -6493772333226108, 833517040657526, 220358442413972, 372755769330, -6868535890317968, 664566135678286, 225755365061283, 2858416831817, -7157521071022387, 490751075721118, 228448778179969, 5269379888994, -7358818790936382, 314165232382833, 228452763163332, 7578988059119, -7471566924126326, 136899005473070, 225812296327790, 9762203913194, -7495942755766923, -38984324020262, 220602211106001, 11795872177577, -7433143529741523, -211472022825831, 212925832011491, 13658956252499, -7285355515665663, -378624356972050, 202913301681642, 15332746247078, -7055712145579987, -538595822537854, 190719625501870, 16801036599608, -6748241887867917, -689654930258378, 176522461172680, 18050271736292, -6367806633571872, -830202339184137, 160519683075597, 19069658617452, -5920031467125852, -958787157130771, 142926753400869, 19851245422781, -5411226778651180, -1074121249927394, 123973933701590, 20389966031698, -4848303747587006, -1175091427164964, 103903371822367, 20683650356548},
		'{2621464726625032, -1601298142322358, -114277463862052, -54557765512014, 3402192470904109, -1521613693668172, -101035526953527, -52555428834631, 4143075592769200, -1441949887694716, -88125723066021, -50522608463608, 4844167648167600, -1362478337710847, -75562184921028, -48464973598293, 5505606112696863, -1283363101544773, -63357707642890, -46388011318305, 6127608592847788, -1204760640672868, -51523776702445, -44297022280332, 6710469021379336, -1126819797494854, -40070597533593, -42197116997554, 7254553845722606, -1049681790049648, -29007126689070, -40093212685504, 7760298217955961, -973480223457764, -18341104403946, -37990030657633, 8228202194534652, -898341117369665, -8079088437780, -35892094253348, 8658826953596720, -824382948694780, 1773510931025, -33803727280864, 9052791037303526, -751716708882984, 11212394882364, -31729052956814, 9410766626308762, -680445975029133, 20234339123843, -29671993324251, 9733475853085184, -610666994071677, 28837156170190, -27636269130411, 10021687160474126, -542468779358319, 37019656947170, -25625400145358, 10276211711460314, -475933218855185, 44781611831263, -23642705902492, 10497899855813746, -411135194280852, 52123711232903, -21691306841762, 10687637658882664, -348142710452834, 59047525827614, -19774125836360, 10846343497467206, -287017034141629, 65555466535792, -17893890083631, 10974964727353150, -227812841736200, 71650744348225, -16053133340965},
		'{2621464726623828, -1601298142322414, -114277463862073, -54557765512018, 3402192470902937, -1521613693668227, -101035526953548, -52555428834635, 4143075592768060, -1441949887694769, -88125723066041, -50522608463611, 4844167648166494, -1362478337710898, -75562184921047, -48464973598296, 5505606112695792, -1283363101544822, -63357707642909, -46388011318308, 6127608592846752, -1204760640672916, -51523776702463, -44297022280336, 6710469021378337, -1126819797494900, -40070597533610, -42197116997558, 7254553845721645, -1049681790049693, -29007126689086, -40093212685508, 7760298217955038, -973480223457806, -18341104403961, -37990030657636, 8228202194533767, -898341117369706, -8079088437795, -35892094253351, 8658826953595873, -824382948694820, 1773510931011, -33803727280867, 9052791037302716, -751716708883021, 11212394882350, -31729052956816, 9410766626307994, -680445975029168, 20234339123830, -29671993324253, 9733475853084454, -610666994071711, 28837156170178, -27636269130413, 10021687160473434, -542468779358351, 37019656947158, -25625400145361, 10276211711459662, -475933218855215, 44781611831252, -23642705902494, 10497899855813134, -411135194280880, 52123711232892, -21691306841764, 10687637658882086, -348142710452861, 59047525827604, -19774125836362, 10846343497466668, -287017034141654, 65555466535783, -17893890083633, 10974964727352650, -227812841736223, 71650744348217, -16053133340967}};
	localparam logic[63:0] Fbi[0:3][0:79] = '{
		'{7789584925020542, 708887221199158, -206702748225345, -19845819841343, 7393588604643268, 873085743790186, -189441643064671, -21110141804839, 6918639246994867, 1024429359565470, -170276674079435, -22108944360993, 6371556198568730, 1161381434685642, -149461551191332, -22835111110926, 5759879607888508, 1282597644249564, -127264837936302, -23284800600437, 5091771080218742, 1386938313763277, -103966594132111, -23457435961284, 4375908801885497, 1473478185138040, -79854941677750, -23355656937657, 3621378440744956, 1541513537288885, -55222594523002, -22985235482842, 2837561156357778, 1590566623196748, -30363393574268, -22354956512906, 2034020064558232, 1620387416998140, -5568886563156, -21476465781011, 1220386496487038, 1630952695911008, 18875008286193, -20364087183631, 406247372102465, 1622462512239921, 42691217575166, -19034612125145, -398965026813756, 1595334139989243, 65614571842042, -17507063846684, -1186079648425665, 1550193608429831, 87394675671855, -15802439866300, -1946288454422587, 1487864961015521, 107798558746626, -13943435878179, -2671242297735851, 1409357402058381, 126613080816752, -11954154617209, -3353139883456778, 1315850515302490, 143647066875003, -9859803310541, -3984808899006887, 1208677757771555, 158733152334642, -7686383409257, -4559778505553668, 1089308448825112, 171729321708043, -5460376320793, -5072342496187033, 959328488094488, 182520128106280, -3208428846785},
		'{-7789584925020678, -708887221199165, 206702748225342, 19845819841342, -7393588604643451, -873085743790196, 189441643064668, 21110141804838, -6918639246995094, -1024429359565484, 170276674079431, 22108944360992, -6371556198568998, -1161381434685658, 149461551191327, 22835111110925, -5759879607888814, -1282597644249583, 127264837936296, 23284800600436, -5091771080219080, -1386938313763298, 103966594132105, 23457435961283, -4375908801885863, -1473478185138064, 79854941677743, 23355656937656, -3621378440745346, -1541513537288910, 55222594522994, 22985235482840, -2837561156358186, -1590566623196775, 30363393574260, 22354956512905, -2034020064558654, -1620387416998168, 5568886563148, 21476465781009, -1220386496487468, -1630952695911038, -18875008286202, 20364087183629, -406247372102900, -1622462512239951, -42691217575174, 19034612125143, 398965026813322, -1595334139989273, -65614571842050, 17507063846682, 1186079648425238, -1550193608429861, -87394675671863, 15802439866299, 1946288454422172, -1487864961015550, -107798558746634, 13943435878177, 2671242297735452, -1409357402058410, -126613080816760, 11954154617207, 3353139883456400, -1315850515302518, -143647066875011, 9859803310540, 3984808899006532, -1208677757771581, -158733152334649, 7686383409256, 4559778505553342, -1089308448825137, -171729321708049, 5460376320792, 5072342496186738, -959328488094511, -182520128106285, 3208428846784},
		'{-20410122023596984, -1087203619517777, -261581401330405, -19688353631198, -19855845437227768, -1129165953014674, -260549776479662, -21497800075813, -19281639300793944, -1166937977762846, -258996978016206, -23185429430581, -18689575854732616, -1200612237457261, -256948048973282, -24752655664962, -18081679793730520, -1230286297560720, -254428064696757, -26201094598827, -17459925861202104, -1256062325165291, -251462077212791, -27532552007075, -16826236651983674, -1278046676369314, -248075061960339, -28749011807856, -16182480619338714, -1296349491750649, -244291866905447, -29852624356494, -15530470282089826, -1311084300475151, -240137164048391, -30845694866052, -14871960627433400, -1322367633538259, -235635403329143, -31730671974348, -14208647704754270, -1330318646597064, -230810768931151, -32510136476076, -13542167405539158, -1335058752810478, -225687137978284, -33186790237559, -12874094424288384, -1336711266066034, -220288041614798, -33763445310536, -12205941395145922, -1335401054933668, -214636628453457, -34243013260277, -11539158198806890, -1331254207649389, -208755630372409, -34628494722203, -10875131434119388, -1324397708395326, -202667330637182, -34922969200132, -10215184048673250, -1314959125107046, -196393534320064, -35129585118164, -9560575122561506, -1303066309004502, -189955540985356, -35251550137213, -8912499799410572, -1288847106009427, -183374119605357, -35292121746123, -8272089358702066, -1272429080179444, -176669485668604, -35254598136332},
		'{20410122023597112, 1087203619517783, 261581401330408, 19688353631199, 19855845437227944, 1129165953014683, 260549776479665, 21497800075814, 19281639300794168, 1166937977762856, 258996978016210, 23185429430582, 18689575854732880, 1200612237457274, 256948048973287, 24752655664963, 18081679793730820, 1230286297560734, 254428064696763, 26201094598828, 17459925861202444, 1256062325165307, 251462077212797, 27532552007076, 16826236651984046, 1278046676369332, 248075061960346, 28749011807857, 16182480619339120, 1296349491750668, 244291866905454, 29852624356495, 15530470282090264, 1311084300475172, 240137164048399, 30845694866053, 14871960627433864, 1322367633538281, 235635403329152, 31730671974350, 14208647704754760, 1330318646597088, 230810768931160, 32510136476078, 13542167405539672, 1335058752810502, 225687137978293, 33186790237561, 12874094424288920, 1336711266066060, 220288041614808, 33763445310538, 12205941395146478, 1335401054933694, 214636628453467, 34243013260279, 11539158198807466, 1331254207649416, 208755630372419, 34628494722205, 10875131434119980, 1324397708395354, 202667330637193, 34922969200134, 10215184048673856, 1314959125107074, 196393534320075, 35129585118166, 9560575122562122, 1303066309004531, 189955540985367, 35251550137215, 8912499799411199, 1288847106009456, 183374119605368, 35292121746125, 8272089358702702, 1272429080179473, 176669485668615, 35254598136334}};
	localparam logic[63:0] hf[0:1999] = {7033096503296, -32897980416, -10967230464, 63928604, 7000245665792, -98394423296, -10337267712, 188110032, 6934845456384, -162997501952, -9086782464, 301512896, 6837488844800, -226124627968, -7233756672, 397524544, 6709056110592, -287210536960, -4804252672, 470098240, 6550703833088, -345713672192, -1831931776, 513814560, 6363853881344, -401122131968, 1642511488, 523933696, 6150172966912, -452959338496, 5571985920, 496438560, 5911558488064, -500788854784, 9903706112, 428068320, 5650113888256, -544219168768, 14579948544, 316342016, 5368126111744, -582907527168, 19538849792, 159572240, 5068042010624, -616563212288, 24715249664, -43130884, 4752438460416, -644950327296, 30041542656, -291865696, 4423997194240, -667889827840, 35448557568, -585954240, 4085474918400, -685260537856, 40866439168, -923966848, 3739673690112, -697000263680, 46225510400, -1303755136, 3389412343808, -703105531904, 51457126400, -1722493184, 3037497131008, -703630671872, 56494514176, -2176726784, 2686692360192, -698686832640, 61273546752, -2662427904, 2339693658112, -688439820288, 65733513216, -3175056896, 1999099920384, -673107279872, 69817778176, -3709628672, 1667389456384, -652956008448, 73474457600, -4260784384, 1346895216640, -628297957376, 76656959488, -4822863872, 1039784017920, -599486234624, 79324479488, -5389984768, 748036685824, -566910648320, 81442447360, -5956117504, 473431015424, -530992660480, 82982838272, -6515166720, 217527091200, -492180406272, 83924451328, -7061048320, -18344486912, -450943287296, 84253073408, -7587765248, -233092038656, -407766368256, 83961561088, -8089484800, -425869180928, -363144806400, 83049857024, -8560607232, -596078428160, -317578280960, 81524924416, -8995835904, -743372095488, -271565209600, 79400542208, -9390236672, -867650306048, -225597456384, 76697108480, -9739302912, -969056190464, -180154810368, 73441320960, -10038998016, -1047968874496, -135700045824, 69665783808, -10285808640, -1104993583104, -92673966080, 65408569344, -10476781568, -1140949254144, -51490967552, 60712722432, -10609551360, -1156854972416, -12534914048, 55625695232, -10682369024, -1153913061376, 23844581376, 50198769664, -10694119424, -1133491388416, 57335398400, 44486422528, -10644324352, -1097103966208, 87665672192, 38545653760, -10533150720, -1046390308864, 114606071808, 32435316736, -10361399296, -983093477376, 137971515392, 26215440384, -10130492416, -909037731840, 157622370304, 19946518528, -9842454528, -826105724928, 173465124864, 13688829952, -9499883520, -736215171072, 185452544000, 7501764608, -9105917952, -641296105472, 193583169536, 1443165440, -8664196096, -543267749888, 197900484608, -4431298048, -8178812416, -444016885760, 198491455488, -10068722688, -7654265856, -345376227328, 195484614656, -15419525120, -7095408640, -249104269312, 189047783424, -20437946368, -6507388928, -156866412544, 179385237504, -25082505216, -5895589888, -70217392128, 166734675968, -29316399104, -5265568768, 9414508544, 151363747840, -33107843072, -4622995968, 80741564416, 133566259200, -36430344192, -3973589248, 142628683776, 113658347520, -39262916608, -3323052544, 194103558144, 91974221824, -41590218752, -2677014272, 234364616704, 68861943808, -43402641408, -2040966400, 262786842624, 44679032832, -44696309760, -1420208256, 278925475840, 19788113920, -45473042432, -819790720, 282517438464, -5447470592, -45740224512, -244465792, 273480531968, -30667960320, -45510623232, 301360416, 251910750208, -55521345536, -44802162688, 813669824, 218077265920, -79667380224, -43637624832, 1288869760, 172415664128, -102781378560, -42044309504, 1723824640, 115519225856, -124557795328, -40053633024, 2115882240, 48128520192, -144713433088, -37700722688, 2462894336, -28880474112, -162990424064, -35023921152, 2763230464, -114509742080, -179158859776, -32064319488, 3015787008, -207653748736, -193018920960, -28865234944, 3219988736, -307115032576, -204402835456, -25471664128, 3375784960, -411620442112, -213176172544, -21929756672, 3483641344, -519838269440, -219238973440, -18286260224, 3544522240, -630395568128, -222526259200, -14587981824, 3559872512, -741895634944, -223008227328, -10881244160, 3531590144, -852935704576, -220690022400, -7211374080, 3461996544, -962124054528, -215611097088, -3622200320, 3353801728, -1068097273856, -207844130816, -155578656, 3210066176, -1169536057344, -197493669888, 3149049344, 3034159104, -1265181130752, -184694308864, 6255063040, 2829713920, -1353847668736, -169608675328, 9129030656, 2600581376, -1434438467584, -152425005056, 11741032448, 2350781696, -1505956593664, -133354577920, 14064936960, 2084455552, -1567515475968, -112628752384, 16078633984, 1805813376, -1618349129728, -90496016384, 17764208640, 1519086592, -1657819234304, -67218747392, 19108071424, 1228478592, -1685421162496, -43069902848, 20101029888, 938116672, -1700789092352, -18329671680, 20738314240, 652006464, -1703698104320, 6717959680, 21019545600, 373988160, -1694065885184, 31788576768, 20948656128, 107695488, -1671951417344, 56600698880, 20533766144, -143481952, -1637553012736, 80879017984, 19787003904, -376432992, -1591204642816, 104357543936, 18724286464, -588355264, -1533370171392, 126782562304, 17365071872, -776781440, -1464636669952, 147915423744, 15732052992, -939601280, -1385706160128, 167535099904, 13850836992, -1075078784, -1297386569728, 185440518144, 11749591040, -1181864704, -1200580722688, 201452535808, 9458661376, -1259004928, -1096275197952, 215415816192, 7010174464, -1305943424, -985527877632, 227200188416, 4437632000, -1322520576, -869455364096, 236701794304, 1775485824, -1308967168, -749219348480, 243843940352, -941283776, -1265894400, -626012913664, 248577572864, -3677590016, -1194278144, -501046935552, 250881425408, -6398656512, -1095440768, -375535730688, 250761838592, -9070423040, -971028672, -250683834368, 248252301312, -11659934720, -822986240, -127672295424, 243412647936, -14135713792, -653526912, -7645917696, 236328009728, -16468104192, -465101920, 108299083776, 227107389440, -18629595136, -260366176, 219126661120, 215882104832, -20595109888, -42143052, 323871637504, 202803920896, -22342254592, 186612704, 421649350656, 188043018240, -23851552768, 422852640, 511664455680, 171785748480, -25106614272, 663472896, 593218240512, 154232242176, -26094284800, 905352320, 665715081216, 135593918464, -26804754432, 1145390336, 728667193344, 116090904576, -27231608832, 1380543744, 781698727936, 95949373440, -27371864064, 1607862400, 824547606528, 75398856704, -27225939968, 1824522752, 857067028480, 54669598720, -26797602816, 2027859968, 879224750080, 33989888000, -26093875200, 2215397376, 891101773824, 13583513600, -25124898816, 2384873216, 892889333760, -6332733440, -23903772672, 2534263552, 884884701184, -25551407104, -22446352384, 2661804288, 867486269440, -43876618240, -20771020800, 2766007296, 841186934784, -61126078464, -18898444288, 2845674240, 806566887424, -77132947456, -16851289088, 2899907328, 764285681664, -91747483648, -14653930496, 2928114688, 715073060864, -104838455296, -12332148736, 2930013696, 659719585792, -116294311936, -9912799232, 2905629696, 599066345472, -126024146944, -7423496704, 2855291904, 533994668032, -133958361088, -4892274176, 2779624704, 465415241728, -140049088512, -2347257600, 2679536640, 394257203200, -144270393344, 183660272, 2556206336, 321457225728, -146618138624, 2673139712, 2411064576, 247948623872, -147109675008, 5094700032, 2245774336, 174650785792, -145783259136, 7423012352, 2062207744, 102458908672, -142697250816, 9634170880, 1862423296, 32234213376, -137929080832, 11705949184, 1648637312, -35205341184, -131574038528, 13618027520, 1423197824, -99093577728, -123743797248, 15352196096, 1188554880, -158723964928, -114564939776, 16892532736, 947231424, -213456617472, -104177123328, 18225549312, 701792896, -262724354048, -92731334656, 19340306432, 454817568, -306037915648, -80387866624, 20228497408, 208866800, -342990127104, -67314339840, 20884506624, -33544018, -373259010048, -53683642368, 21305427968, -269973504, -396609880064, -39671808000, 21491048448, -498081024, -412896460800, -25455941632, 21443817472, -715651776, -422060851200, -11212149760, 21168769024, -920620160, -424132542464, 2886491648, 20673421312, -1111091072, -419226353664, 16671883264, 19967651840, -1285358592, -407539548160, 29982767104, 19063545856, -1441922816, -389347966976, 42666471424, 17975222272, -1579503232, -365001244672, 54580543488, 16718628864, -1697049984, -334917435392, 65594208256, 15311344640, -1793752448, -299576754176, 75589697536, 13772339200, -1869043840, -259514777600, 84463378432, 12121732096, -1922604416, -215315218432, 92126724096, 10380551168, -1954360704, -167602061312, 98507071488, 8570467840, -1964482176, -117031575552, 103548190720, 6713540096, -1953375744, -64283930624, 107210645504, 4831954432, -1921676416, -10054776832, 109471981568, 2947766016, -1870237312, 44953247744, 110326685696, 1082651264, -1800114816, 100038934528, 109785948160, -742337920, -1712554752, 154510770176, 107877253120, -2507003392, -1608973312, 207694921728, 104643788800, -4192218624, -1490939392, 258942943232, 100143644672, -5780130304, -1360152832, 307638960128, 94448910336, -7254341120, -1218423808, 353206403072, 87644585984, -8600073216, -1067649472, 395114184704, 79827378176, -9804311552, -909791232, 432882253824, 71104356352, -10855919616, -746850816, 466086363136, 61591547904, -11745739776, -580847104, 494362230784, 51412426752, -12466658304, -413792224, 517408784384, 40696356864, -13013656576, -247669072, 534990848000, 29576974336, -13383830528, -84408840, 546940780544, 18190557184, -13576387584, 74130096, 553159360512, 6674405888, -13592614912, 226182256, 553615949824, -4834780672, -13435834368, 370093632, 548347740160, -16202491904, -13111324672, 504338656, 537458442240, -27297931264, -12626223104, 627535488, 521115828224, -37995479040, -11989416960, 738459264, 499548880896, -48176078848, -11211404288, 836053504, 473044221952, -57728499712, -10304146432, 919438912, 441941950464, -66550517760, -9280902144, 987920768, 406630694912, -74549952512, -8156052992, 1040993088, 367542566912, -81645584384, -6944914944, 1078341504, 325147328512, -87767891968, -5663543808, 1099843200, 279946461184, -92859727872, -4328539136, 1105564672, 232466825216, -96876699648, -2956838144, 1095757824, 183254220800, -99787579392, -1565513600, 1070853440, 132866760704, -101574352896, -171574784, 1031453312, 81868210176, -102232301568, 1208231424, 978319616, 30821447680, -101769781248, 2557609472, 912363520, -19718068224, -100207943680, 3860898560, 834631680, -69208547328, -97580294144, 5103242240, 746291840, -117127929856, -93932068864, 6270749696, 648616768, -162979545088, -89319563264, 7350639104, 542967744, -206297481216, -83809280000, 8331369472, 430777056, -246651437056, -77476986880, 9202753536, 313529888, -283651080192, -70406725632, 9956050944, 192746128, -316949954560, -62689660928, 10584052736, 69961976, -346248708096, -54422949888, 11081128960, -53288364, -371297878016, -45708509184, 11443279872, -175490560, -391899774976, -36651757568, 11668144128, -295167552, -407910121472, -27360344064, 11755006976, -410896192, -419238739968, -17942872064, 11704777728, -521323040, -425849716736, -8507630592, 11519951872, -625179008, -427760877568, 838650880, 11204558848, -721292672, -425042903040, 9992007680, 10764085248, -808602688, -417817427968, 18852395008, 10205391872, -886167872, -406254944256, 27324768256, 9536608256, -953176704, -390571982848, 35320111104, 8767017984, -1008954368, -371027836928, 42756349952, 7906931200, -1052968640, -347921055744, 49559191552, 6967550976, -1084833536, -321585086464, 55662837760, 5960825344, -1104311424, -292384145408, 61010624512, 4899297280, -1111313664, -260708253696, 65555509248, 3795950592, -1105899136, -226968616960, 69260451840, 2664050688, -1088270976, -191592300544, 72098676736, 1516986752, -1058772032, -155017199616, 74053804032, 368114528, -1017878592, -117686788096, 75119886336, -769398208, -966192896, -80044908544, 75301273600, -1882721152, -904433792, -42530721792, 74612400128, -2959504384, -833426688, -5573702144, 73077473280, -3988013824, -754092160, 30411114496, 70729965568, -4957257216, -667433984, 65027657728, 67612160000, -5857098752, -574525888, 97903050752, 63774429184, -6678363136, -476498048, 128691486720, 59274575872, -7412924928, -374523168, 157077749760, 54177009664, -8053787136, -269802144, 182780313600, 48551907328, -8595142656, -163549664, 205553975296, 42474287104, -9032420352, -56980000, 225192067072, 36023083008, -9362321408, 48707084, 241528176640, 29280149504, -9582834688, 152339968, 254437326848, 22329272320, -9693236224, 252788304, 263836680192, 15255162880, -9694081024, 348975392, 269685833728, 8142476288, -9587174400, 439889728, 271986458624, 1074818560, -9375527936, 524595744, 270781579264, -5866192896, -9063308288, 602243328, 266154344448, -12601840640, -8655766528, 672076160, 258226323456, -19057170432, -8159164928, 733439296, 247155507200, -25161789440, -7580680704, 785784512, 233133752320, -30850611200, -6928315392, 828675456, 216383995904, -36064505856, -6210783744, 861790464, 197157126144, -40750891008, -5437403136, 884924608, 175728607232, -44864233472, -4617976320, 897990272, 152394776576, -48366440448, -3762670080, 901015872, 127469125632, -51227189248, -2881891584, 894144000, 101278294016, -53424144384, -1986164096, 877627648, 74158080000, -54943068160, -1086004096, 851825792, 46449369088, -55777853440, -191799792, 817197120, 18494062592, -55930470400, 686306496, 774293504, -9368892416, -55410786304, 1538531200, 723751744, -36807413760, -54236319744, 2355556864, 666285184, -63500029952, -52431921152, 3128631040, 602673856, -89139437568, -50029350912, 3849658368, 533754816, -113435836416, -47066787840, 4511283200, 460411168, -136120008704, -43588292608, 5106960896, 383561312, -156946137088, -39643185152, 5631021568, 304147840, -175694184448, -35285385216, 6078718976, 223126112, -192172146688, -30572709888, 6446269952, 141453168, -206217691136, -25566150656, 6730883584, 60076656, -217699647488, -20329084928, 6930774016, -20075964, -226518974464, -14926526464, 7045166592, -98107728, -232609366016, -9424327680, 7074288128, -173161984, -235937497088, -3888407296, 7019345920, -244431584, -236502859776, 1616015232, 6882502144, -311167360, -234337206272, 7025165824, 6666826240, -372685728, -229503696896, 12277432320, 6376248320, -428375552, -222095589376, 17314041856, 6015498752, -477703744, -212234715136, 22079696896, 5590036992, -520220320, -200069513216, 26523152384, 5105980416, -555562048, -185772982272, 30597754880, 4570017280, -583455104, -169540141056, 34261897216, 3989324800, -603716864, -151585505280, 37479415808, 3371473408, -616256256, -132140228608, 40219930624, 2724335104, -621073344, -111449161728, 42459090944, 2055986048, -618257728, -89767772160, 44178755584, 1374610176, -607985920, -67359031296, 45367111680, 688401792, -590518080, -44490215424, 46018699264, 5471468, -566193024, -21429762048, 46134370304, -666247424, -535423520, 1555883136, 45721169920, -1319086976, -498689888, 24205301760, 44792164352, -1945729536, -456533408, 46265061376, 43366166528, -2539286272, -409548928, 67492519936, 41467457536, -3093369600, -358377120, 87658446848, 39125377024, -3602159872, -303696256, 106549485568, 36373929984, -4060461568, -246213632, 123970330624, 33251299328, -4463754240, -186656976, 139745705984, 29799337984, -4808232448, -125765560, 153722093568, 26063024128, -5090839552, -64281496, 165769084928, 22089889792, -5309289472, -2941044, 175780577280, 17929424896, -5462078464, 57533836, 183675584512, 13632480256, -5548493312, 116443600, 189398745088, 9250644992, -5568603136, 173118880, 192920535040, 4835645952, -5523246592, 226927712, 194237251584, 438742560, -5414009344, 277282272, 193370537984, -3889856000, -5243192832, 323644960, 190366760960, -8101555712, -5013775360, 365533728, 185296093184, -12149912576, -4729367040, 402526848, 178251268096, -15991135232, -4394157056, 434266688, 169346187264, -19584544768, -4012854528, 460462816, 158714167296, -22892994560, -3590626816, 480894272, 146506186752, -25883242496, -3133030656, 495411008, 132888772608, -28526272512, -2645941760, 503934304, 118041862144, -30797553664, -2135481216, 506456576, 102156492800, -32677253120, -1607940736, 503040352, 85432393728, -34150387712, -1069706688, 493816192, 68075581440, -35206914048, -527184576, 478980192, 50295820288, -35841761280, 13275691, 458790528, 32304191488, -36054810624, 545452224, 433563520, 14310600704, -35850821632, 1063321216, 403668896, -3478606336, -35239272448, 1561123456, 369524608, -20862973952, -34234189824, 2033426688, 331591296, -37650149376, -32853913600, 2475182848, 290366144, -53657956352, -31120795648, 2881780480, 246376544, -68716351488, -29060892672, 3249091072, 200173424, -82669150208, -26703589376, 3573507840, 152324528, -95375622144, -24081211392, 3851980032, 103407576, -106711851008, -21228597248, 4082038528, 54003312, -116571865088, -18182653952, 4261814272, 4688806, -124868567040, -14981902336, 4390051328, -43969216, -131534446592, -11665993728, 4466109440, -91420760, -136521965568, -8275239936, 4489962496, -137138640, -139803836416, -4850135552, 4462188544, -180624272, -141372964864, -1430882688, 4383951872, -221412864, -141242171392, 1943064960, 4256981760, -259078384, -139443732480, 5233448448, 4083541248, -293237696, -136028684288, 8403623936, 3866393344, -323554464, -131065856000, 11418961920, 3608760064, -349742080, -124640845824, 14247211008, 3314277632, -371566368, -116854710272, 16858833920, 2986947328, -388847200, -107822514176, 19227299840, 2631084288, -401459936, -97671798784, 21329344512, 2251260672, -409335712, -86540869632, 23145181184, 1852249216, -412461504, -74577018880, 24658677760, 1438965504, -410879232, -61934665728, 25857468416, 1016407424, -404684448, -48773451776, 26733047808, 589596736, -394024256, -35256303616, 27280797696, 163520480, -379094880, -21547479040, 27499972608, -256926192, -360138432, -7810651136, 27393648640, -666995136, -337439520, 5792974336, 26968619008, -1062137472, -311321088, 19106494464, 26235260928, -1438052992, -282140192, 31979048960, 25207339008, -1790736000, -250283168, 44267466752, 23901808640, -2116516096, -216160832, 55837798400, 22338547712, -2412095488, -180203184, 66566709248, 20540094464, -2674580480, -142854208, 76342730752, 18531325952, -2901509120, -104566496, 85067358208, 16339141632, -3090871296, -65795828, 92655960064, 13992113152, -3241124864, -26995910, 99038543872, 11520123904, -3351205888, 11386859, 104160296960, 8954007552, -3420532224, 48918428, 107981996032, 6325167616, -3449003264, 85181896, 110480179200, 3665207808, -3436992256, 119782032, 111647170560, 1005561408, -3385333760, 152349504, 111490867200, -1622868352, -3295307008, 182544688, 110034436096, -4190059008, -3168613632, 210061120, 107315757056, -6667201024, -3007350016, 234628432, 103386734592, -9027011584, -2813977088, 256014944, 98312503296, -11244024832, -2591285760, 274029632, 92170379264, -13294855168, -2342358784, 288523648, 85048827904, -15158435840, -2070530560, 299391392, 77046226944, -16816222208, -1779343616, 306570976, 68269547520, -18252363776, -1472505088, 310044160, 58832982016, -19453847552, -1153840384, 309835904, 48856506368, -20410593280, -827246976, 306013216, 38464389120, -21115523072, -496648352, 298683904, 27783663616, -21564604416, -165947968, 287994368, 16942639104, -21756829696, 161015488, 274127456, 6069367296, -21694183424, 480511552, 257299680, -4709823488, -21381576704, 788959168, 237758064, -15271768064, -20826730496, 1082965888, 215776896, -25497839616, -20040044544, 1359363712, 191653968, -35275247616, -19034429440, 1615242112, 165706880, -44498239488, -17825124352, 1847977472, 138268864, -53069225984, -16429464576, 2055258368, 109684824, -60899762176, -14866663424, 2235107584, 80307000, -67911417856, -13157547008, 2385898752, 50490892, -74036527104, -11324291072, 2506369792, 20591002, -79218802688, -9390139392, 2595631104, -9043209, -83413778432, -7379118592, 2653169920, -38071296, -86589120512, -5315746304, 2678849792, -66165620, -88724840448, -3224739072, 2672905216, -93014920, -89813286912, -1130721792, 2635934208, -118327656, -89859039232, 942053824, 2568883456, -141835040, -88878645248, 2969985280, 2473032960, -163293760, -86900252672, 4930381312, 2349974784, -182488384, -83963068416, 6801708544, 2201590016, -199233408, -80116711424, 8563822592, 2030020992, -213374832, -75420508160, 10198177792, 1837643904, -224791472, -69942599680, 11688014848, 1627035520, -233395808, -63759036416, 13018524672, 1400941312, -239134400, -56952745984, 14176988160, 1162240128, -241988000, -49612476416, 15152887808, 913908864, -241971088, -41831669760, 15937992704, 658986304, -239131280, -33707284480, 16526415872, 400536864, -233548080, -25338644480, 16914642944, 141614768, -225331520, -16826230784, 17101535232, -114771248, -214620368, -8270504960, 17088299008, -365691968, -201579968, 229250672, 16878435328, -608330368, -186399968, 8576060928, 16477662208, -840012160, -169291648, 16676343808, 15893807104, -1058234624, -150485136, 24440932352, 15136688128, -1260692480, -130226448, 31786033152, 14217958400, -1445301760, -108774312, 38634110976, 13150946304, -1610219392, -86397032, 44914671616, 11950475264, -1753861248, -63369172, 50564964352, 10632657920, -1874915968, -39968276, 55530573824, 9214700544, -1972355584, -16471616, 59765919744, 7714673664, -2045442560, 6847026, 63234625536, 6151298560, -2093733376, 29720462, 65909788672, 4543711744, -2117079296, 51891092, 67774132224, 2911243008, -2115622528, 73113720, 68820041728, 1273183616, -2089790208, 93158192, 69049499648, -351433280, -2040284416, 111811808, 68473896960, -1944049536, -1968069376, 128881496, 67113725952, -3486789120, -1874356352, 144195728, 64998219776, -4962652672, -1760584960, 157606112, 62164844544, -6355700736, -1628403200, 168988784, 58658750464, -7651218944, -1479644416, 178245392, 54532087808, -8835868672, -1316303360, 185303792, 49843318784, -9897820160, -1140510208, 190118496, 44656418816, -10826858496, -954503680, 192670752, 39040032768, -11614480384, -760603392, 192968256, 33066635264, -12253963264, -561181504, 191044672, 26811590656, -12740410368, -358634592, 186958800, 20352258048, -13070778368, -155355344, 180793488, 13767048192, -13243881472, 46295076, 172654240, 7134508032, -13260374016, 244013680, 162667648, 532402080, -13122712576, 435581472, 150979568, -5963171840, -12835095552, 618887680, 137753088, -12278635520, -12403388416, 791952384, 123166384, -18343737344, -11835023360, 952947136, 107410400, -24092315648, -11138892800, 1100213760, 90686408, -29462990848, -10325217280, 1232280576, 73203528, -34399793152, -9405405184, 1347876480, 55176152, -38852730880, -8391904768, 1445942016, 36821416, -42778251264, -7298036736, 1525638272, 18356602, -46139658240, -6137830912, 1586352896, -3364, -48907403264, -4925849088, 1627703296, -18048354, -51059314688, -3677007104, 1649537408, -35575396, -52580737024, -2406398464, 1651931392, -52390896, -53464559616, -1129114624, 1635185152, -68312728, -53711183872, 139928944, 1599814784, -83172152, -53328396288, 1386162304, 1546543488, -96815528, -52331134976, 2595524096, 1476289152, -109105848, -50741219328, 3754616064, 1390150784, -119924056, -48586973184, 4850846208, 1289392896, -129170104, -45902774272, 5872562688, 1175427840, -136763808, -42728583168, 6809170432, 1049796992, -142645424, -39109353472, 7651239424, 914150976, -146776032, -35094458368, 8390590464, 770228544, -149137584, -30737025024, 9020372992, 619834944, -149732832, -26093264896, 9535118336, 464820192, -148584864, -21221765120, 9930782720, 307056544, -145736576, -16182777856, 10204768256, 148416656, -141249808, -11037487104, 10355931136, -9248055, -135204288, -5847291392, 10384567296, -164128624, -127696448, -673083584, 10292387840, -314478656, -118838032, 4425443328, 10082473984, -458633504, -108754496, 9390467072, 9759219712, -595028224, -97583376, 14166675456, 9328256000, -722214016, -85472480, 18701864960, 8796367872, -838872960, -72578000, 22947489792, 8171397632, -943831040, -59062548, 26859171840, 7462130688, -1036069504, -45093212, 30397132800, 6678184448, -1114734080, -30839494, 33526589440, 5829879808, -1179141760, -16471352, 36218060800, 4928109056, -1228786048, -2157196, 38447636480, 3984203008, -1263340160, 11938022, 40197140480, 3009790464, -1282657280, 25654662, 41454268416, 2016659712, -1286769408, 38840152, 42212614144, 1016618176, -1275884288, 51350640, 42471653376, 21356334, -1250379776, 63052516, 42236645376, -957685888, -1210796416, 73823768, 41518489600, -1909447296, -1157828864, 83555224, 40333484032, -2823367424, -1092315392, 92151592, 38703067136, -3689500160, -1015224960, 99532312, 36653469696, -4498618368, -927644736, 105632264, 34215340032, -5242309120, -830765056, 110402272, 31423309824, -5913057792, -725863872, 113809368, 28315527168, -6504319488, -614290688, 115836928, 24933158912, -7010576896, -497449664, 116484592, 21319860224, -7427391488, -376782464, 115767992, 17521235968, -7751432704, -253750912, 113718288, 13584269312, -7980498432, -129819680, 110381560, 9556759552, -8113524224, -6439408, 105818040, 5486758400, -8150574080, 114969968, 100101136, 1422006400, -8092821504, 233035072, 93316416, -2590614528, -7942518272, 346444256, 85560352, -6505608704, -7702948864, 453961664, 76939064, -10279368704, -7378376192, 554440448, 67566928, -13870651392, -6973975552, 646834304, 57565096, -17241012224, -6495759872, 730208128, 47059976, -20355205120, -5950494720, 803746816, 36181704, -23181537280, -5345609216, 866762944, 25062552, -25692176384, -4689098240, 918702144, 13835381, -27863408640, -3989420544, 959147840, 2632072, -29675841536, -3255392000, 987823232, -8417969, -31114557440, -2496078848, 1004592512, -19189274, -32169211904, -1720688896, 1009460096, -29561700, -32834078720, -938460864, 1002568000, -39421732, -33108035584, -158558640, 984192000, -48663680, -32994498560, 610034432, 954736192, -57190776};
	localparam logic[63:0] hb[0:1999] = {7033096503296, 32897980416, -10967230464, -63928604, 7000245665792, 98394423296, -10337267712, -188110032, 6934845456384, 162997501952, -9086782464, -301512896, 6837488844800, 226124627968, -7233756672, -397524544, 6709056110592, 287210536960, -4804252672, -470098240, 6550703833088, 345713672192, -1831931776, -513814560, 6363853881344, 401122131968, 1642511488, -523933696, 6150172966912, 452959338496, 5571985920, -496438560, 5911558488064, 500788854784, 9903706112, -428068320, 5650113888256, 544219168768, 14579948544, -316342016, 5368126111744, 582907527168, 19538849792, -159572240, 5068042010624, 616563212288, 24715249664, 43130884, 4752438460416, 644950327296, 30041542656, 291865696, 4423997194240, 667889827840, 35448557568, 585954240, 4085474918400, 685260537856, 40866439168, 923966848, 3739673690112, 697000263680, 46225510400, 1303755136, 3389412343808, 703105531904, 51457126400, 1722493184, 3037497131008, 703630671872, 56494514176, 2176726784, 2686692360192, 698686832640, 61273546752, 2662427904, 2339693658112, 688439820288, 65733513216, 3175056896, 1999099920384, 673107279872, 69817778176, 3709628672, 1667389456384, 652956008448, 73474457600, 4260784384, 1346895216640, 628297957376, 76656959488, 4822863872, 1039784017920, 599486234624, 79324479488, 5389984768, 748036685824, 566910648320, 81442447360, 5956117504, 473431015424, 530992660480, 82982838272, 6515166720, 217527091200, 492180406272, 83924451328, 7061048320, -18344486912, 450943287296, 84253073408, 7587765248, -233092038656, 407766368256, 83961561088, 8089484800, -425869180928, 363144806400, 83049857024, 8560607232, -596078428160, 317578280960, 81524924416, 8995835904, -743372095488, 271565209600, 79400542208, 9390236672, -867650306048, 225597456384, 76697108480, 9739302912, -969056190464, 180154810368, 73441320960, 10038998016, -1047968874496, 135700045824, 69665783808, 10285808640, -1104993583104, 92673966080, 65408569344, 10476781568, -1140949254144, 51490967552, 60712722432, 10609551360, -1156854972416, 12534914048, 55625695232, 10682369024, -1153913061376, -23844581376, 50198769664, 10694119424, -1133491388416, -57335398400, 44486422528, 10644324352, -1097103966208, -87665672192, 38545653760, 10533150720, -1046390308864, -114606071808, 32435316736, 10361399296, -983093477376, -137971515392, 26215440384, 10130492416, -909037731840, -157622370304, 19946518528, 9842454528, -826105724928, -173465124864, 13688829952, 9499883520, -736215171072, -185452544000, 7501764608, 9105917952, -641296105472, -193583169536, 1443165440, 8664196096, -543267749888, -197900484608, -4431298048, 8178812416, -444016885760, -198491455488, -10068722688, 7654265856, -345376227328, -195484614656, -15419525120, 7095408640, -249104269312, -189047783424, -20437946368, 6507388928, -156866412544, -179385237504, -25082505216, 5895589888, -70217392128, -166734675968, -29316399104, 5265568768, 9414508544, -151363747840, -33107843072, 4622995968, 80741564416, -133566259200, -36430344192, 3973589248, 142628683776, -113658347520, -39262916608, 3323052544, 194103558144, -91974221824, -41590218752, 2677014272, 234364616704, -68861943808, -43402641408, 2040966400, 262786842624, -44679032832, -44696309760, 1420208256, 278925475840, -19788113920, -45473042432, 819790720, 282517438464, 5447470592, -45740224512, 244465792, 273480531968, 30667960320, -45510623232, -301360416, 251910750208, 55521345536, -44802162688, -813669824, 218077265920, 79667380224, -43637624832, -1288869760, 172415664128, 102781378560, -42044309504, -1723824640, 115519225856, 124557795328, -40053633024, -2115882240, 48128520192, 144713433088, -37700722688, -2462894336, -28880474112, 162990424064, -35023921152, -2763230464, -114509742080, 179158859776, -32064319488, -3015787008, -207653748736, 193018920960, -28865234944, -3219988736, -307115032576, 204402835456, -25471664128, -3375784960, -411620442112, 213176172544, -21929756672, -3483641344, -519838269440, 219238973440, -18286260224, -3544522240, -630395568128, 222526259200, -14587981824, -3559872512, -741895634944, 223008227328, -10881244160, -3531590144, -852935704576, 220690022400, -7211374080, -3461996544, -962124054528, 215611097088, -3622200320, -3353801728, -1068097273856, 207844130816, -155578656, -3210066176, -1169536057344, 197493669888, 3149049344, -3034159104, -1265181130752, 184694308864, 6255063040, -2829713920, -1353847668736, 169608675328, 9129030656, -2600581376, -1434438467584, 152425005056, 11741032448, -2350781696, -1505956593664, 133354577920, 14064936960, -2084455552, -1567515475968, 112628752384, 16078633984, -1805813376, -1618349129728, 90496016384, 17764208640, -1519086592, -1657819234304, 67218747392, 19108071424, -1228478592, -1685421162496, 43069902848, 20101029888, -938116672, -1700789092352, 18329671680, 20738314240, -652006464, -1703698104320, -6717959680, 21019545600, -373988160, -1694065885184, -31788576768, 20948656128, -107695488, -1671951417344, -56600698880, 20533766144, 143481952, -1637553012736, -80879017984, 19787003904, 376432992, -1591204642816, -104357543936, 18724286464, 588355264, -1533370171392, -126782562304, 17365071872, 776781440, -1464636669952, -147915423744, 15732052992, 939601280, -1385706160128, -167535099904, 13850836992, 1075078784, -1297386569728, -185440518144, 11749591040, 1181864704, -1200580722688, -201452535808, 9458661376, 1259004928, -1096275197952, -215415816192, 7010174464, 1305943424, -985527877632, -227200188416, 4437632000, 1322520576, -869455364096, -236701794304, 1775485824, 1308967168, -749219348480, -243843940352, -941283776, 1265894400, -626012913664, -248577572864, -3677590016, 1194278144, -501046935552, -250881425408, -6398656512, 1095440768, -375535730688, -250761838592, -9070423040, 971028672, -250683834368, -248252301312, -11659934720, 822986240, -127672295424, -243412647936, -14135713792, 653526912, -7645917696, -236328009728, -16468104192, 465101920, 108299083776, -227107389440, -18629595136, 260366176, 219126661120, -215882104832, -20595109888, 42143052, 323871637504, -202803920896, -22342254592, -186612704, 421649350656, -188043018240, -23851552768, -422852640, 511664455680, -171785748480, -25106614272, -663472896, 593218240512, -154232242176, -26094284800, -905352320, 665715081216, -135593918464, -26804754432, -1145390336, 728667193344, -116090904576, -27231608832, -1380543744, 781698727936, -95949373440, -27371864064, -1607862400, 824547606528, -75398856704, -27225939968, -1824522752, 857067028480, -54669598720, -26797602816, -2027859968, 879224750080, -33989888000, -26093875200, -2215397376, 891101773824, -13583513600, -25124898816, -2384873216, 892889333760, 6332733440, -23903772672, -2534263552, 884884701184, 25551407104, -22446352384, -2661804288, 867486269440, 43876618240, -20771020800, -2766007296, 841186934784, 61126078464, -18898444288, -2845674240, 806566887424, 77132947456, -16851289088, -2899907328, 764285681664, 91747483648, -14653930496, -2928114688, 715073060864, 104838455296, -12332148736, -2930013696, 659719585792, 116294311936, -9912799232, -2905629696, 599066345472, 126024146944, -7423496704, -2855291904, 533994668032, 133958361088, -4892274176, -2779624704, 465415241728, 140049088512, -2347257600, -2679536640, 394257203200, 144270393344, 183660272, -2556206336, 321457225728, 146618138624, 2673139712, -2411064576, 247948623872, 147109675008, 5094700032, -2245774336, 174650785792, 145783259136, 7423012352, -2062207744, 102458908672, 142697250816, 9634170880, -1862423296, 32234213376, 137929080832, 11705949184, -1648637312, -35205341184, 131574038528, 13618027520, -1423197824, -99093577728, 123743797248, 15352196096, -1188554880, -158723964928, 114564939776, 16892532736, -947231424, -213456617472, 104177123328, 18225549312, -701792896, -262724354048, 92731334656, 19340306432, -454817568, -306037915648, 80387866624, 20228497408, -208866800, -342990127104, 67314339840, 20884506624, 33544018, -373259010048, 53683642368, 21305427968, 269973504, -396609880064, 39671808000, 21491048448, 498081024, -412896460800, 25455941632, 21443817472, 715651776, -422060851200, 11212149760, 21168769024, 920620160, -424132542464, -2886491648, 20673421312, 1111091072, -419226353664, -16671883264, 19967651840, 1285358592, -407539548160, -29982767104, 19063545856, 1441922816, -389347966976, -42666471424, 17975222272, 1579503232, -365001244672, -54580543488, 16718628864, 1697049984, -334917435392, -65594208256, 15311344640, 1793752448, -299576754176, -75589697536, 13772339200, 1869043840, -259514777600, -84463378432, 12121732096, 1922604416, -215315218432, -92126724096, 10380551168, 1954360704, -167602061312, -98507071488, 8570467840, 1964482176, -117031575552, -103548190720, 6713540096, 1953375744, -64283930624, -107210645504, 4831954432, 1921676416, -10054776832, -109471981568, 2947766016, 1870237312, 44953247744, -110326685696, 1082651264, 1800114816, 100038934528, -109785948160, -742337920, 1712554752, 154510770176, -107877253120, -2507003392, 1608973312, 207694921728, -104643788800, -4192218624, 1490939392, 258942943232, -100143644672, -5780130304, 1360152832, 307638960128, -94448910336, -7254341120, 1218423808, 353206403072, -87644585984, -8600073216, 1067649472, 395114184704, -79827378176, -9804311552, 909791232, 432882253824, -71104356352, -10855919616, 746850816, 466086363136, -61591547904, -11745739776, 580847104, 494362230784, -51412426752, -12466658304, 413792224, 517408784384, -40696356864, -13013656576, 247669072, 534990848000, -29576974336, -13383830528, 84408840, 546940780544, -18190557184, -13576387584, -74130096, 553159360512, -6674405888, -13592614912, -226182256, 553615949824, 4834780672, -13435834368, -370093632, 548347740160, 16202491904, -13111324672, -504338656, 537458442240, 27297931264, -12626223104, -627535488, 521115828224, 37995479040, -11989416960, -738459264, 499548880896, 48176078848, -11211404288, -836053504, 473044221952, 57728499712, -10304146432, -919438912, 441941950464, 66550517760, -9280902144, -987920768, 406630694912, 74549952512, -8156052992, -1040993088, 367542566912, 81645584384, -6944914944, -1078341504, 325147328512, 87767891968, -5663543808, -1099843200, 279946461184, 92859727872, -4328539136, -1105564672, 232466825216, 96876699648, -2956838144, -1095757824, 183254220800, 99787579392, -1565513600, -1070853440, 132866760704, 101574352896, -171574784, -1031453312, 81868210176, 102232301568, 1208231424, -978319616, 30821447680, 101769781248, 2557609472, -912363520, -19718068224, 100207943680, 3860898560, -834631680, -69208547328, 97580294144, 5103242240, -746291840, -117127929856, 93932068864, 6270749696, -648616768, -162979545088, 89319563264, 7350639104, -542967744, -206297481216, 83809280000, 8331369472, -430777056, -246651437056, 77476986880, 9202753536, -313529888, -283651080192, 70406725632, 9956050944, -192746128, -316949954560, 62689660928, 10584052736, -69961976, -346248708096, 54422949888, 11081128960, 53288364, -371297878016, 45708509184, 11443279872, 175490560, -391899774976, 36651757568, 11668144128, 295167552, -407910121472, 27360344064, 11755006976, 410896192, -419238739968, 17942872064, 11704777728, 521323040, -425849716736, 8507630592, 11519951872, 625179008, -427760877568, -838650880, 11204558848, 721292672, -425042903040, -9992007680, 10764085248, 808602688, -417817427968, -18852395008, 10205391872, 886167872, -406254944256, -27324768256, 9536608256, 953176704, -390571982848, -35320111104, 8767017984, 1008954368, -371027836928, -42756349952, 7906931200, 1052968640, -347921055744, -49559191552, 6967550976, 1084833536, -321585086464, -55662837760, 5960825344, 1104311424, -292384145408, -61010624512, 4899297280, 1111313664, -260708253696, -65555509248, 3795950592, 1105899136, -226968616960, -69260451840, 2664050688, 1088270976, -191592300544, -72098676736, 1516986752, 1058772032, -155017199616, -74053804032, 368114528, 1017878592, -117686788096, -75119886336, -769398208, 966192896, -80044908544, -75301273600, -1882721152, 904433792, -42530721792, -74612400128, -2959504384, 833426688, -5573702144, -73077473280, -3988013824, 754092160, 30411114496, -70729965568, -4957257216, 667433984, 65027657728, -67612160000, -5857098752, 574525888, 97903050752, -63774429184, -6678363136, 476498048, 128691486720, -59274575872, -7412924928, 374523168, 157077749760, -54177009664, -8053787136, 269802144, 182780313600, -48551907328, -8595142656, 163549664, 205553975296, -42474287104, -9032420352, 56980000, 225192067072, -36023083008, -9362321408, -48707084, 241528176640, -29280149504, -9582834688, -152339968, 254437326848, -22329272320, -9693236224, -252788304, 263836680192, -15255162880, -9694081024, -348975392, 269685833728, -8142476288, -9587174400, -439889728, 271986458624, -1074818560, -9375527936, -524595744, 270781579264, 5866192896, -9063308288, -602243328, 266154344448, 12601840640, -8655766528, -672076160, 258226323456, 19057170432, -8159164928, -733439296, 247155507200, 25161789440, -7580680704, -785784512, 233133752320, 30850611200, -6928315392, -828675456, 216383995904, 36064505856, -6210783744, -861790464, 197157126144, 40750891008, -5437403136, -884924608, 175728607232, 44864233472, -4617976320, -897990272, 152394776576, 48366440448, -3762670080, -901015872, 127469125632, 51227189248, -2881891584, -894144000, 101278294016, 53424144384, -1986164096, -877627648, 74158080000, 54943068160, -1086004096, -851825792, 46449369088, 55777853440, -191799792, -817197120, 18494062592, 55930470400, 686306496, -774293504, -9368892416, 55410786304, 1538531200, -723751744, -36807413760, 54236319744, 2355556864, -666285184, -63500029952, 52431921152, 3128631040, -602673856, -89139437568, 50029350912, 3849658368, -533754816, -113435836416, 47066787840, 4511283200, -460411168, -136120008704, 43588292608, 5106960896, -383561312, -156946137088, 39643185152, 5631021568, -304147840, -175694184448, 35285385216, 6078718976, -223126112, -192172146688, 30572709888, 6446269952, -141453168, -206217691136, 25566150656, 6730883584, -60076656, -217699647488, 20329084928, 6930774016, 20075964, -226518974464, 14926526464, 7045166592, 98107728, -232609366016, 9424327680, 7074288128, 173161984, -235937497088, 3888407296, 7019345920, 244431584, -236502859776, -1616015232, 6882502144, 311167360, -234337206272, -7025165824, 6666826240, 372685728, -229503696896, -12277432320, 6376248320, 428375552, -222095589376, -17314041856, 6015498752, 477703744, -212234715136, -22079696896, 5590036992, 520220320, -200069513216, -26523152384, 5105980416, 555562048, -185772982272, -30597754880, 4570017280, 583455104, -169540141056, -34261897216, 3989324800, 603716864, -151585505280, -37479415808, 3371473408, 616256256, -132140228608, -40219930624, 2724335104, 621073344, -111449161728, -42459090944, 2055986048, 618257728, -89767772160, -44178755584, 1374610176, 607985920, -67359031296, -45367111680, 688401792, 590518080, -44490215424, -46018699264, 5471468, 566193024, -21429762048, -46134370304, -666247424, 535423520, 1555883136, -45721169920, -1319086976, 498689888, 24205301760, -44792164352, -1945729536, 456533408, 46265061376, -43366166528, -2539286272, 409548928, 67492519936, -41467457536, -3093369600, 358377120, 87658446848, -39125377024, -3602159872, 303696256, 106549485568, -36373929984, -4060461568, 246213632, 123970330624, -33251299328, -4463754240, 186656976, 139745705984, -29799337984, -4808232448, 125765560, 153722093568, -26063024128, -5090839552, 64281496, 165769084928, -22089889792, -5309289472, 2941044, 175780577280, -17929424896, -5462078464, -57533836, 183675584512, -13632480256, -5548493312, -116443600, 189398745088, -9250644992, -5568603136, -173118880, 192920535040, -4835645952, -5523246592, -226927712, 194237251584, -438742560, -5414009344, -277282272, 193370537984, 3889856000, -5243192832, -323644960, 190366760960, 8101555712, -5013775360, -365533728, 185296093184, 12149912576, -4729367040, -402526848, 178251268096, 15991135232, -4394157056, -434266688, 169346187264, 19584544768, -4012854528, -460462816, 158714167296, 22892994560, -3590626816, -480894272, 146506186752, 25883242496, -3133030656, -495411008, 132888772608, 28526272512, -2645941760, -503934304, 118041862144, 30797553664, -2135481216, -506456576, 102156492800, 32677253120, -1607940736, -503040352, 85432393728, 34150387712, -1069706688, -493816192, 68075581440, 35206914048, -527184576, -478980192, 50295820288, 35841761280, 13275691, -458790528, 32304191488, 36054810624, 545452224, -433563520, 14310600704, 35850821632, 1063321216, -403668896, -3478606336, 35239272448, 1561123456, -369524608, -20862973952, 34234189824, 2033426688, -331591296, -37650149376, 32853913600, 2475182848, -290366144, -53657956352, 31120795648, 2881780480, -246376544, -68716351488, 29060892672, 3249091072, -200173424, -82669150208, 26703589376, 3573507840, -152324528, -95375622144, 24081211392, 3851980032, -103407576, -106711851008, 21228597248, 4082038528, -54003312, -116571865088, 18182653952, 4261814272, -4688806, -124868567040, 14981902336, 4390051328, 43969216, -131534446592, 11665993728, 4466109440, 91420760, -136521965568, 8275239936, 4489962496, 137138640, -139803836416, 4850135552, 4462188544, 180624272, -141372964864, 1430882688, 4383951872, 221412864, -141242171392, -1943064960, 4256981760, 259078384, -139443732480, -5233448448, 4083541248, 293237696, -136028684288, -8403623936, 3866393344, 323554464, -131065856000, -11418961920, 3608760064, 349742080, -124640845824, -14247211008, 3314277632, 371566368, -116854710272, -16858833920, 2986947328, 388847200, -107822514176, -19227299840, 2631084288, 401459936, -97671798784, -21329344512, 2251260672, 409335712, -86540869632, -23145181184, 1852249216, 412461504, -74577018880, -24658677760, 1438965504, 410879232, -61934665728, -25857468416, 1016407424, 404684448, -48773451776, -26733047808, 589596736, 394024256, -35256303616, -27280797696, 163520480, 379094880, -21547479040, -27499972608, -256926192, 360138432, -7810651136, -27393648640, -666995136, 337439520, 5792974336, -26968619008, -1062137472, 311321088, 19106494464, -26235260928, -1438052992, 282140192, 31979048960, -25207339008, -1790736000, 250283168, 44267466752, -23901808640, -2116516096, 216160832, 55837798400, -22338547712, -2412095488, 180203184, 66566709248, -20540094464, -2674580480, 142854208, 76342730752, -18531325952, -2901509120, 104566496, 85067358208, -16339141632, -3090871296, 65795828, 92655960064, -13992113152, -3241124864, 26995910, 99038543872, -11520123904, -3351205888, -11386859, 104160296960, -8954007552, -3420532224, -48918428, 107981996032, -6325167616, -3449003264, -85181896, 110480179200, -3665207808, -3436992256, -119782032, 111647170560, -1005561408, -3385333760, -152349504, 111490867200, 1622868352, -3295307008, -182544688, 110034436096, 4190059008, -3168613632, -210061120, 107315757056, 6667201024, -3007350016, -234628432, 103386734592, 9027011584, -2813977088, -256014944, 98312503296, 11244024832, -2591285760, -274029632, 92170379264, 13294855168, -2342358784, -288523648, 85048827904, 15158435840, -2070530560, -299391392, 77046226944, 16816222208, -1779343616, -306570976, 68269547520, 18252363776, -1472505088, -310044160, 58832982016, 19453847552, -1153840384, -309835904, 48856506368, 20410593280, -827246976, -306013216, 38464389120, 21115523072, -496648352, -298683904, 27783663616, 21564604416, -165947968, -287994368, 16942639104, 21756829696, 161015488, -274127456, 6069367296, 21694183424, 480511552, -257299680, -4709823488, 21381576704, 788959168, -237758064, -15271768064, 20826730496, 1082965888, -215776896, -25497839616, 20040044544, 1359363712, -191653968, -35275247616, 19034429440, 1615242112, -165706880, -44498239488, 17825124352, 1847977472, -138268864, -53069225984, 16429464576, 2055258368, -109684824, -60899762176, 14866663424, 2235107584, -80307000, -67911417856, 13157547008, 2385898752, -50490892, -74036527104, 11324291072, 2506369792, -20591002, -79218802688, 9390139392, 2595631104, 9043209, -83413778432, 7379118592, 2653169920, 38071296, -86589120512, 5315746304, 2678849792, 66165620, -88724840448, 3224739072, 2672905216, 93014920, -89813286912, 1130721792, 2635934208, 118327656, -89859039232, -942053824, 2568883456, 141835040, -88878645248, -2969985280, 2473032960, 163293760, -86900252672, -4930381312, 2349974784, 182488384, -83963068416, -6801708544, 2201590016, 199233408, -80116711424, -8563822592, 2030020992, 213374832, -75420508160, -10198177792, 1837643904, 224791472, -69942599680, -11688014848, 1627035520, 233395808, -63759036416, -13018524672, 1400941312, 239134400, -56952745984, -14176988160, 1162240128, 241988000, -49612476416, -15152887808, 913908864, 241971088, -41831669760, -15937992704, 658986304, 239131280, -33707284480, -16526415872, 400536864, 233548080, -25338644480, -16914642944, 141614768, 225331520, -16826230784, -17101535232, -114771248, 214620368, -8270504960, -17088299008, -365691968, 201579968, 229250672, -16878435328, -608330368, 186399968, 8576060928, -16477662208, -840012160, 169291648, 16676343808, -15893807104, -1058234624, 150485136, 24440932352, -15136688128, -1260692480, 130226448, 31786033152, -14217958400, -1445301760, 108774312, 38634110976, -13150946304, -1610219392, 86397032, 44914671616, -11950475264, -1753861248, 63369172, 50564964352, -10632657920, -1874915968, 39968276, 55530573824, -9214700544, -1972355584, 16471616, 59765919744, -7714673664, -2045442560, -6847026, 63234625536, -6151298560, -2093733376, -29720462, 65909788672, -4543711744, -2117079296, -51891092, 67774132224, -2911243008, -2115622528, -73113720, 68820041728, -1273183616, -2089790208, -93158192, 69049499648, 351433280, -2040284416, -111811808, 68473896960, 1944049536, -1968069376, -128881496, 67113725952, 3486789120, -1874356352, -144195728, 64998219776, 4962652672, -1760584960, -157606112, 62164844544, 6355700736, -1628403200, -168988784, 58658750464, 7651218944, -1479644416, -178245392, 54532087808, 8835868672, -1316303360, -185303792, 49843318784, 9897820160, -1140510208, -190118496, 44656418816, 10826858496, -954503680, -192670752, 39040032768, 11614480384, -760603392, -192968256, 33066635264, 12253963264, -561181504, -191044672, 26811590656, 12740410368, -358634592, -186958800, 20352258048, 13070778368, -155355344, -180793488, 13767048192, 13243881472, 46295076, -172654240, 7134508032, 13260374016, 244013680, -162667648, 532402080, 13122712576, 435581472, -150979568, -5963171840, 12835095552, 618887680, -137753088, -12278635520, 12403388416, 791952384, -123166384, -18343737344, 11835023360, 952947136, -107410400, -24092315648, 11138892800, 1100213760, -90686408, -29462990848, 10325217280, 1232280576, -73203528, -34399793152, 9405405184, 1347876480, -55176152, -38852730880, 8391904768, 1445942016, -36821416, -42778251264, 7298036736, 1525638272, -18356602, -46139658240, 6137830912, 1586352896, 3364, -48907403264, 4925849088, 1627703296, 18048354, -51059314688, 3677007104, 1649537408, 35575396, -52580737024, 2406398464, 1651931392, 52390896, -53464559616, 1129114624, 1635185152, 68312728, -53711183872, -139928944, 1599814784, 83172152, -53328396288, -1386162304, 1546543488, 96815528, -52331134976, -2595524096, 1476289152, 109105848, -50741219328, -3754616064, 1390150784, 119924056, -48586973184, -4850846208, 1289392896, 129170104, -45902774272, -5872562688, 1175427840, 136763808, -42728583168, -6809170432, 1049796992, 142645424, -39109353472, -7651239424, 914150976, 146776032, -35094458368, -8390590464, 770228544, 149137584, -30737025024, -9020372992, 619834944, 149732832, -26093264896, -9535118336, 464820192, 148584864, -21221765120, -9930782720, 307056544, 145736576, -16182777856, -10204768256, 148416656, 141249808, -11037487104, -10355931136, -9248055, 135204288, -5847291392, -10384567296, -164128624, 127696448, -673083584, -10292387840, -314478656, 118838032, 4425443328, -10082473984, -458633504, 108754496, 9390467072, -9759219712, -595028224, 97583376, 14166675456, -9328256000, -722214016, 85472480, 18701864960, -8796367872, -838872960, 72578000, 22947489792, -8171397632, -943831040, 59062548, 26859171840, -7462130688, -1036069504, 45093212, 30397132800, -6678184448, -1114734080, 30839494, 33526589440, -5829879808, -1179141760, 16471352, 36218060800, -4928109056, -1228786048, 2157196, 38447636480, -3984203008, -1263340160, -11938022, 40197140480, -3009790464, -1282657280, -25654662, 41454268416, -2016659712, -1286769408, -38840152, 42212614144, -1016618176, -1275884288, -51350640, 42471653376, -21356334, -1250379776, -63052516, 42236645376, 957685888, -1210796416, -73823768, 41518489600, 1909447296, -1157828864, -83555224, 40333484032, 2823367424, -1092315392, -92151592, 38703067136, 3689500160, -1015224960, -99532312, 36653469696, 4498618368, -927644736, -105632264, 34215340032, 5242309120, -830765056, -110402272, 31423309824, 5913057792, -725863872, -113809368, 28315527168, 6504319488, -614290688, -115836928, 24933158912, 7010576896, -497449664, -116484592, 21319860224, 7427391488, -376782464, -115767992, 17521235968, 7751432704, -253750912, -113718288, 13584269312, 7980498432, -129819680, -110381560, 9556759552, 8113524224, -6439408, -105818040, 5486758400, 8150574080, 114969968, -100101136, 1422006400, 8092821504, 233035072, -93316416, -2590614528, 7942518272, 346444256, -85560352, -6505608704, 7702948864, 453961664, -76939064, -10279368704, 7378376192, 554440448, -67566928, -13870651392, 6973975552, 646834304, -57565096, -17241012224, 6495759872, 730208128, -47059976, -20355205120, 5950494720, 803746816, -36181704, -23181537280, 5345609216, 866762944, -25062552, -25692176384, 4689098240, 918702144, -13835381, -27863408640, 3989420544, 959147840, -2632072, -29675841536, 3255392000, 987823232, 8417969, -31114557440, 2496078848, 1004592512, 19189274, -32169211904, 1720688896, 1009460096, 29561700, -32834078720, 938460864, 1002568000, 39421732, -33108035584, 158558640, 984192000, 48663680, -32994498560, -610034432, 954736192, 57190776};
endpackage
`endif
