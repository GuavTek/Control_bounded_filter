`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam N = 4;
	localparam M = 4;
	localparam real Lfr[0:3] = {0.9909936, 0.9909936, 0.9798975, 0.9798975};
	localparam real Lfi[0:3] = {0.04006346, -0.04006346, 0.016101336, -0.016101336};
	localparam real Lbr[0:3] = {0.9909936, 0.9909936, 0.9798975, 0.9798975};
	localparam real Lbi[0:3] = {0.04006346, -0.04006346, 0.016101336, -0.016101336};
	localparam real Wfr[0:3] = {-6.379518e-06, -6.379518e-06, -1.8966227e-06, -1.8966227e-06};
	localparam real Wfi[0:3] = {-2.512436e-07, 2.512436e-07, -3.6578447e-06, 3.6578447e-06};
	localparam real Wbr[0:3] = {6.379518e-06, 6.379518e-06, 1.8966227e-06, 1.8966227e-06};
	localparam real Wbi[0:3] = {2.512436e-07, -2.512436e-07, 3.6578447e-06, -3.6578447e-06};
	localparam real Ffr[0:3][0:99] = '{
		'{-315.39786, -25.729626, 2.391748, -0.02091026, -327.88712, -24.224422, 2.4033616, -0.026568063, -339.61957, -22.702948, 2.4107327, -0.032088693, -350.58783, -21.168032, 2.413919, -0.037465084, -360.78583, -19.62248, 2.4129825, -0.042690527, -370.20898, -18.069077, 2.4079926, -0.04775867, -378.85406, -16.510567, 2.399024, -0.052663535, -386.71915, -14.949662, 2.3861566, -0.05739952, -393.80377, -13.389033, 2.3694756, -0.061961398, -400.10867, -11.831307, 2.3490715, -0.06634431, -405.636, -10.279063, 2.3250399, -0.0705438, -410.38907, -8.73483, 2.2974799, -0.074555784, -414.37256, -7.2010803, 2.2664957, -0.07837655, -417.5923, -5.6802287, 2.2321959, -0.08200277, -420.05533, -4.1746297, 2.1946921, -0.08543151, -421.76984, -2.6865723, 2.1541, -0.088660225, -422.7452, -1.2182797, 2.1105382, -0.091686726, -422.9918, 0.22809494, 2.0641289, -0.09450921, -422.5211, 1.6504707, 2.0149968, -0.09712625, -421.34564, 3.046841, 1.9632692, -0.09953679, -419.4789, 4.415276, 1.9090756, -0.101740144, -416.93533, 5.753924, 1.8525478, -0.10373596, -413.73026, 7.061014, 1.7938192, -0.10552428, -409.87985, 8.334858, 1.7330246, -0.107105464, -405.40118, 9.57385, 1.6703004, -0.10848024},
		'{-315.39786, -25.729626, 2.391748, -0.02091026, -327.88712, -24.224422, 2.4033616, -0.026568063, -339.61957, -22.702948, 2.4107327, -0.032088693, -350.58783, -21.168032, 2.413919, -0.037465084, -360.78583, -19.62248, 2.4129825, -0.042690527, -370.20898, -18.069077, 2.4079926, -0.04775867, -378.85406, -16.510567, 2.399024, -0.052663535, -386.71915, -14.949662, 2.3861566, -0.05739952, -393.80377, -13.389033, 2.3694756, -0.061961398, -400.10867, -11.831307, 2.3490715, -0.06634431, -405.636, -10.279063, 2.3250399, -0.0705438, -410.38907, -8.73483, 2.2974799, -0.074555784, -414.37256, -7.2010803, 2.2664957, -0.07837655, -417.5923, -5.6802287, 2.2321959, -0.08200277, -420.05533, -4.1746297, 2.1946921, -0.08543151, -421.76984, -2.6865723, 2.1541, -0.088660225, -422.7452, -1.2182797, 2.1105382, -0.091686726, -422.9918, 0.22809494, 2.0641289, -0.09450921, -422.5211, 1.6504707, 2.0149968, -0.09712625, -421.34564, 3.046841, 1.9632692, -0.09953679, -419.4789, 4.415276, 1.9090756, -0.101740144, -416.93533, 5.753924, 1.8525478, -0.10373596, -413.73026, 7.061014, 1.7938192, -0.10552428, -409.87985, 8.334858, 1.7330246, -0.107105464, -405.40118, 9.57385, 1.6703004, -0.10848024},
		'{-313.9008, -25.617615, 2.3192613, -0.26458496, -326.34842, -24.179775, 2.2132473, -0.25634763, -338.08737, -22.782751, 2.1099567, -0.24826594, -349.13785, -21.425854, 2.009351, -0.24033912, -359.51978, -20.108398, 1.9113904, -0.23256631, -369.25272, -18.829697, 1.8160353, -0.22494659, -378.35583, -17.589067, 1.7232461, -0.21747893, -386.848, -16.385826, 1.6329827, -0.21016228, -394.74777, -15.219293, 1.5452054, -0.20299554, -402.0733, -14.08879, 1.4598737, -0.19597752, -408.84244, -12.993643, 1.3769478, -0.189107, -415.07272, -11.933181, 1.2963876, -0.1823827, -420.78128, -10.906735, 1.2181528, -0.17580332, -425.98502, -9.913642, 1.1422035, -0.16936746, -430.70038, -8.95324, 1.0684996, -0.16307375, -434.94357, -8.024876, 0.9970013, -0.1569207, -438.73047, -7.1278963, 0.9276688, -0.15090688, -442.0766, -6.2616568, 0.8604624, -0.14503074, -444.99716, -5.425516, 0.79534274, -0.13929075, -447.50702, -4.618839, 0.73227036, -0.13368532, -449.6208, -3.8409946, 0.67120624, -0.12821287, -451.35272, -3.0913596, 0.6121114, -0.12287174, -452.71674, -2.3693159, 0.5549472, -0.11766031, -453.72653, -1.6742512, 0.49967527, -0.112576894, -454.3954, -1.0055599, 0.44625738, -0.1076198},
		'{-313.9008, -25.617615, 2.3192613, -0.26458496, -326.34842, -24.179775, 2.2132473, -0.25634763, -338.08737, -22.782751, 2.1099567, -0.24826594, -349.13785, -21.425854, 2.009351, -0.24033912, -359.51978, -20.108398, 1.9113904, -0.23256631, -369.25272, -18.829697, 1.8160353, -0.22494659, -378.35583, -17.589067, 1.7232461, -0.21747893, -386.848, -16.385826, 1.6329827, -0.21016228, -394.74777, -15.219293, 1.5452054, -0.20299554, -402.0733, -14.08879, 1.4598737, -0.19597752, -408.84244, -12.993643, 1.3769478, -0.189107, -415.07272, -11.933181, 1.2963876, -0.1823827, -420.78128, -10.906735, 1.2181528, -0.17580332, -425.98502, -9.913642, 1.1422035, -0.16936746, -430.70038, -8.95324, 1.0684996, -0.16307375, -434.94357, -8.024876, 0.9970013, -0.1569207, -438.73047, -7.1278963, 0.9276688, -0.15090688, -442.0766, -6.2616568, 0.8604624, -0.14503074, -444.99716, -5.425516, 0.79534274, -0.13929075, -447.50702, -4.618839, 0.73227036, -0.13368532, -449.6208, -3.8409946, 0.67120624, -0.12821287, -451.35272, -3.0913596, 0.6121114, -0.12287174, -452.71674, -2.3693159, 0.5549472, -0.11766031, -453.72653, -1.6742512, 0.49967527, -0.112576894, -454.3954, -1.0055599, 0.44625738, -0.1076198}};
	localparam real Ffi[0:3][0:99] = '{
		'{382.63885, -31.786383, -0.82754797, 0.1459217, 366.55676, -32.530922, -0.7242731, 0.14376976, 350.1191, -33.20845, -0.621463, 0.1414105, 333.35947, -33.81892, -0.5192836, 0.13885131, 316.31137, -34.3624, -0.4178968, 0.1360998, 299.0082, -34.839066, -0.31746066, 0.1331637, 281.48337, -35.249203, -0.21812896, 0.130051, 263.77005, -35.593204, -0.12005121, 0.12676983, 245.90112, -35.871574, -0.023372298, 0.12332847, 227.9093, -36.08491, 0.07176759, 0.119735345, 209.82693, -36.23392, 0.16523317, 0.11599898, 191.68597, -36.3194, 0.25689414, 0.11212802, 173.51797, -36.342243, 0.34662545, 0.10813119, 155.354, -36.303432, 0.43430728, 0.10401729, 137.22464, -36.204037, 0.5198252, 0.099795155, 119.159874, -36.045223, 0.60307044, 0.095473684, 101.18912, -35.82822, 0.6839397, 0.09106178, 83.34113, -35.554344, 0.76233536, 0.086568356, 65.64402, -35.22499, 0.8381656, 0.08200232, 48.12515, -34.841618, 0.9113445, 0.077372566, 30.811152, -34.405754, 0.981792, 0.07268793, 13.72788, -33.918995, 1.0494338, 0.067957215, -3.0996308, -33.382984, 1.1142017, 0.06318915, -19.64718, -32.799435, 1.1760334, 0.058392372, -35.891434, -32.17011, 1.2348726, 0.053575456},
		'{-382.63885, 31.786383, 0.82754797, -0.1459217, -366.55676, 32.530922, 0.7242731, -0.14376976, -350.1191, 33.20845, 0.621463, -0.1414105, -333.35947, 33.81892, 0.5192836, -0.13885131, -316.31137, 34.3624, 0.4178968, -0.1360998, -299.0082, 34.839066, 0.31746066, -0.1331637, -281.48337, 35.249203, 0.21812896, -0.130051, -263.77005, 35.593204, 0.12005121, -0.12676983, -245.90112, 35.871574, 0.023372298, -0.12332847, -227.9093, 36.08491, -0.07176759, -0.119735345, -209.82693, 36.23392, -0.16523317, -0.11599898, -191.68597, 36.3194, -0.25689414, -0.11212802, -173.51797, 36.342243, -0.34662545, -0.10813119, -155.354, 36.303432, -0.43430728, -0.10401729, -137.22464, 36.204037, -0.5198252, -0.099795155, -119.159874, 36.045223, -0.60307044, -0.095473684, -101.18912, 35.82822, -0.6839397, -0.09106178, -83.34113, 35.554344, -0.76233536, -0.086568356, -65.64402, 35.22499, -0.8381656, -0.08200232, -48.12515, 34.841618, -0.9113445, -0.077372566, -30.811152, 34.405754, -0.981792, -0.07268793, -13.72788, 33.918995, -1.0494338, -0.067957215, 3.0996308, 33.382984, -1.1142017, -0.06318915, 19.64718, 32.799435, -1.1760334, -0.058392372, 35.891434, 32.17011, -1.2348726, -0.053575456},
		'{1164.9854, -57.3158, 3.6885912, -0.18126035, 1136.5121, -56.576088, 3.6517847, -0.18187673, 1108.4106, -55.828094, 3.6140108, -0.1823481, 1080.6852, -55.072643, 3.5753334, -0.18267986, 1053.3391, -54.31053, 3.5358136, -0.18287732, 1026.3756, -53.542526, 3.4955108, -0.18294565, 999.7974, -52.76937, 3.4544828, -0.18288992, 973.607, -51.991783, 3.4127858, -0.18271509, 947.8063, -51.21045, 3.3704734, -0.18242595, 922.39703, -50.426044, 3.3275983, -0.18202724, 897.3806, -49.639202, 3.2842112, -0.18152353, 872.7581, -48.850544, 3.240361, -0.18091933, 848.5303, -48.06067, 3.1960952, -0.18021901, 824.6976, -47.27014, 3.1514597, -0.17942682, 801.2602, -46.479515, 3.1064985, -0.17854694, 778.218, -45.68932, 3.0612543, -0.1775834, 755.5707, -44.900063, 3.0157685, -0.17654017, 733.3177, -44.11223, 2.9700809, -0.17542107, 711.4581, -43.326283, 2.9242294, -0.17422986, 689.991, -42.542675, 2.878251, -0.17297018, 668.91504, -41.76183, 2.8321817, -0.17164555, 648.22864, -40.984158, 2.786055, -0.17025945, 627.93024, -40.21005, 2.7399042, -0.1688152, 608.01794, -39.439877, 2.6937606, -0.16731608, 588.4897, -38.673992, 2.6476548, -0.16576526},
		'{-1164.9854, 57.3158, -3.6885912, 0.18126035, -1136.5121, 56.576088, -3.6517847, 0.18187673, -1108.4106, 55.828094, -3.6140108, 0.1823481, -1080.6852, 55.072643, -3.5753334, 0.18267986, -1053.3391, 54.31053, -3.5358136, 0.18287732, -1026.3756, 53.542526, -3.4955108, 0.18294565, -999.7974, 52.76937, -3.4544828, 0.18288992, -973.607, 51.991783, -3.4127858, 0.18271509, -947.8063, 51.21045, -3.3704734, 0.18242595, -922.39703, 50.426044, -3.3275983, 0.18202724, -897.3806, 49.639202, -3.2842112, 0.18152353, -872.7581, 48.850544, -3.240361, 0.18091933, -848.5303, 48.06067, -3.1960952, 0.18021901, -824.6976, 47.27014, -3.1514597, 0.17942682, -801.2602, 46.479515, -3.1064985, 0.17854694, -778.218, 45.68932, -3.0612543, 0.1775834, -755.5707, 44.900063, -3.0157685, 0.17654017, -733.3177, 44.11223, -2.9700809, 0.17542107, -711.4581, 43.326283, -2.9242294, 0.17422986, -689.991, 42.542675, -2.878251, 0.17297018, -668.91504, 41.76183, -2.8321817, 0.17164555, -648.22864, 40.984158, -2.786055, 0.17025945, -627.93024, 40.21005, -2.7399042, 0.1688152, -608.01794, 39.439877, -2.6937606, 0.16731608, -588.4897, 38.673992, -2.6476548, 0.16576526}};
	localparam real Fbr[0:3][0:99] = '{
		'{315.39786, -25.729626, -2.391748, -0.02091026, 327.88712, -24.224422, -2.4033616, -0.026568063, 339.61957, -22.702948, -2.4107327, -0.032088693, 350.58783, -21.168032, -2.413919, -0.037465084, 360.78583, -19.62248, -2.4129825, -0.042690527, 370.20898, -18.069077, -2.4079926, -0.04775867, 378.85406, -16.510567, -2.399024, -0.052663535, 386.71915, -14.949662, -2.3861566, -0.05739952, 393.80377, -13.389033, -2.3694756, -0.061961398, 400.10867, -11.831307, -2.3490715, -0.06634431, 405.636, -10.279063, -2.3250399, -0.0705438, 410.38907, -8.73483, -2.2974799, -0.074555784, 414.37256, -7.2010803, -2.2664957, -0.07837655, 417.5923, -5.6802287, -2.2321959, -0.08200277, 420.05533, -4.1746297, -2.1946921, -0.08543151, 421.76984, -2.6865723, -2.1541, -0.088660225, 422.7452, -1.2182797, -2.1105382, -0.091686726, 422.9918, 0.22809494, -2.0641289, -0.09450921, 422.5211, 1.6504707, -2.0149968, -0.09712625, 421.34564, 3.046841, -1.9632692, -0.09953679, 419.4789, 4.415276, -1.9090756, -0.101740144, 416.93533, 5.753924, -1.8525478, -0.10373596, 413.73026, 7.061014, -1.7938192, -0.10552428, 409.87985, 8.334858, -1.7330246, -0.107105464, 405.40118, 9.57385, -1.6703004, -0.10848024},
		'{315.39786, -25.729626, -2.391748, -0.02091026, 327.88712, -24.224422, -2.4033616, -0.026568063, 339.61957, -22.702948, -2.4107327, -0.032088693, 350.58783, -21.168032, -2.413919, -0.037465084, 360.78583, -19.62248, -2.4129825, -0.042690527, 370.20898, -18.069077, -2.4079926, -0.04775867, 378.85406, -16.510567, -2.399024, -0.052663535, 386.71915, -14.949662, -2.3861566, -0.05739952, 393.80377, -13.389033, -2.3694756, -0.061961398, 400.10867, -11.831307, -2.3490715, -0.06634431, 405.636, -10.279063, -2.3250399, -0.0705438, 410.38907, -8.73483, -2.2974799, -0.074555784, 414.37256, -7.2010803, -2.2664957, -0.07837655, 417.5923, -5.6802287, -2.2321959, -0.08200277, 420.05533, -4.1746297, -2.1946921, -0.08543151, 421.76984, -2.6865723, -2.1541, -0.088660225, 422.7452, -1.2182797, -2.1105382, -0.091686726, 422.9918, 0.22809494, -2.0641289, -0.09450921, 422.5211, 1.6504707, -2.0149968, -0.09712625, 421.34564, 3.046841, -1.9632692, -0.09953679, 419.4789, 4.415276, -1.9090756, -0.101740144, 416.93533, 5.753924, -1.8525478, -0.10373596, 413.73026, 7.061014, -1.7938192, -0.10552428, 409.87985, 8.334858, -1.7330246, -0.107105464, 405.40118, 9.57385, -1.6703004, -0.10848024},
		'{313.9008, -25.617615, -2.3192613, -0.26458496, 326.34842, -24.179775, -2.2132473, -0.25634763, 338.08737, -22.782751, -2.1099567, -0.24826594, 349.13785, -21.425854, -2.009351, -0.24033912, 359.51978, -20.108398, -1.9113904, -0.23256631, 369.25272, -18.829697, -1.8160353, -0.22494659, 378.35583, -17.589067, -1.7232461, -0.21747893, 386.848, -16.385826, -1.6329827, -0.21016228, 394.74777, -15.219293, -1.5452054, -0.20299554, 402.0733, -14.08879, -1.4598737, -0.19597752, 408.84244, -12.993643, -1.3769478, -0.189107, 415.07272, -11.933181, -1.2963876, -0.1823827, 420.78128, -10.906735, -1.2181528, -0.17580332, 425.98502, -9.913642, -1.1422035, -0.16936746, 430.70038, -8.95324, -1.0684996, -0.16307375, 434.94357, -8.024876, -0.9970013, -0.1569207, 438.73047, -7.1278963, -0.9276688, -0.15090688, 442.0766, -6.2616568, -0.8604624, -0.14503074, 444.99716, -5.425516, -0.79534274, -0.13929075, 447.50702, -4.618839, -0.73227036, -0.13368532, 449.6208, -3.8409946, -0.67120624, -0.12821287, 451.35272, -3.0913596, -0.6121114, -0.12287174, 452.71674, -2.3693159, -0.5549472, -0.11766031, 453.72653, -1.6742512, -0.49967527, -0.112576894, 454.3954, -1.0055599, -0.44625738, -0.1076198},
		'{313.9008, -25.617615, -2.3192613, -0.26458496, 326.34842, -24.179775, -2.2132473, -0.25634763, 338.08737, -22.782751, -2.1099567, -0.24826594, 349.13785, -21.425854, -2.009351, -0.24033912, 359.51978, -20.108398, -1.9113904, -0.23256631, 369.25272, -18.829697, -1.8160353, -0.22494659, 378.35583, -17.589067, -1.7232461, -0.21747893, 386.848, -16.385826, -1.6329827, -0.21016228, 394.74777, -15.219293, -1.5452054, -0.20299554, 402.0733, -14.08879, -1.4598737, -0.19597752, 408.84244, -12.993643, -1.3769478, -0.189107, 415.07272, -11.933181, -1.2963876, -0.1823827, 420.78128, -10.906735, -1.2181528, -0.17580332, 425.98502, -9.913642, -1.1422035, -0.16936746, 430.70038, -8.95324, -1.0684996, -0.16307375, 434.94357, -8.024876, -0.9970013, -0.1569207, 438.73047, -7.1278963, -0.9276688, -0.15090688, 442.0766, -6.2616568, -0.8604624, -0.14503074, 444.99716, -5.425516, -0.79534274, -0.13929075, 447.50702, -4.618839, -0.73227036, -0.13368532, 449.6208, -3.8409946, -0.67120624, -0.12821287, 451.35272, -3.0913596, -0.6121114, -0.12287174, 452.71674, -2.3693159, -0.5549472, -0.11766031, 453.72653, -1.6742512, -0.49967527, -0.112576894, 454.3954, -1.0055599, -0.44625738, -0.1076198}};
	localparam real Fbi[0:3][0:99] = '{
		'{-382.63885, -31.786383, 0.82754797, 0.1459217, -366.55676, -32.530922, 0.7242731, 0.14376976, -350.1191, -33.20845, 0.621463, 0.1414105, -333.35947, -33.81892, 0.5192836, 0.13885131, -316.31137, -34.3624, 0.4178968, 0.1360998, -299.0082, -34.839066, 0.31746066, 0.1331637, -281.48337, -35.249203, 0.21812896, 0.130051, -263.77005, -35.593204, 0.12005121, 0.12676983, -245.90112, -35.871574, 0.023372298, 0.12332847, -227.9093, -36.08491, -0.07176759, 0.119735345, -209.82693, -36.23392, -0.16523317, 0.11599898, -191.68597, -36.3194, -0.25689414, 0.11212802, -173.51797, -36.342243, -0.34662545, 0.10813119, -155.354, -36.303432, -0.43430728, 0.10401729, -137.22464, -36.204037, -0.5198252, 0.099795155, -119.159874, -36.045223, -0.60307044, 0.095473684, -101.18912, -35.82822, -0.6839397, 0.09106178, -83.34113, -35.554344, -0.76233536, 0.086568356, -65.64402, -35.22499, -0.8381656, 0.08200232, -48.12515, -34.841618, -0.9113445, 0.077372566, -30.811152, -34.405754, -0.981792, 0.07268793, -13.72788, -33.918995, -1.0494338, 0.067957215, 3.0996308, -33.382984, -1.1142017, 0.06318915, 19.64718, -32.799435, -1.1760334, 0.058392372, 35.891434, -32.17011, -1.2348726, 0.053575456},
		'{382.63885, 31.786383, -0.82754797, -0.1459217, 366.55676, 32.530922, -0.7242731, -0.14376976, 350.1191, 33.20845, -0.621463, -0.1414105, 333.35947, 33.81892, -0.5192836, -0.13885131, 316.31137, 34.3624, -0.4178968, -0.1360998, 299.0082, 34.839066, -0.31746066, -0.1331637, 281.48337, 35.249203, -0.21812896, -0.130051, 263.77005, 35.593204, -0.12005121, -0.12676983, 245.90112, 35.871574, -0.023372298, -0.12332847, 227.9093, 36.08491, 0.07176759, -0.119735345, 209.82693, 36.23392, 0.16523317, -0.11599898, 191.68597, 36.3194, 0.25689414, -0.11212802, 173.51797, 36.342243, 0.34662545, -0.10813119, 155.354, 36.303432, 0.43430728, -0.10401729, 137.22464, 36.204037, 0.5198252, -0.099795155, 119.159874, 36.045223, 0.60307044, -0.095473684, 101.18912, 35.82822, 0.6839397, -0.09106178, 83.34113, 35.554344, 0.76233536, -0.086568356, 65.64402, 35.22499, 0.8381656, -0.08200232, 48.12515, 34.841618, 0.9113445, -0.077372566, 30.811152, 34.405754, 0.981792, -0.07268793, 13.72788, 33.918995, 1.0494338, -0.067957215, -3.0996308, 33.382984, 1.1142017, -0.06318915, -19.64718, 32.799435, 1.1760334, -0.058392372, -35.891434, 32.17011, 1.2348726, -0.053575456},
		'{-1164.9854, -57.3158, -3.6885912, -0.18126035, -1136.5121, -56.576088, -3.6517847, -0.18187673, -1108.4106, -55.828094, -3.6140108, -0.1823481, -1080.6852, -55.072643, -3.5753334, -0.18267986, -1053.3391, -54.31053, -3.5358136, -0.18287732, -1026.3756, -53.542526, -3.4955108, -0.18294565, -999.7974, -52.76937, -3.4544828, -0.18288992, -973.607, -51.991783, -3.4127858, -0.18271509, -947.8063, -51.21045, -3.3704734, -0.18242595, -922.39703, -50.426044, -3.3275983, -0.18202724, -897.3806, -49.639202, -3.2842112, -0.18152353, -872.7581, -48.850544, -3.240361, -0.18091933, -848.5303, -48.06067, -3.1960952, -0.18021901, -824.6976, -47.27014, -3.1514597, -0.17942682, -801.2602, -46.479515, -3.1064985, -0.17854694, -778.218, -45.68932, -3.0612543, -0.1775834, -755.5707, -44.900063, -3.0157685, -0.17654017, -733.3177, -44.11223, -2.9700809, -0.17542107, -711.4581, -43.326283, -2.9242294, -0.17422986, -689.991, -42.542675, -2.878251, -0.17297018, -668.91504, -41.76183, -2.8321817, -0.17164555, -648.22864, -40.984158, -2.786055, -0.17025945, -627.93024, -40.21005, -2.7399042, -0.1688152, -608.01794, -39.439877, -2.6937606, -0.16731608, -588.4897, -38.673992, -2.6476548, -0.16576526},
		'{1164.9854, 57.3158, 3.6885912, 0.18126035, 1136.5121, 56.576088, 3.6517847, 0.18187673, 1108.4106, 55.828094, 3.6140108, 0.1823481, 1080.6852, 55.072643, 3.5753334, 0.18267986, 1053.3391, 54.31053, 3.5358136, 0.18287732, 1026.3756, 53.542526, 3.4955108, 0.18294565, 999.7974, 52.76937, 3.4544828, 0.18288992, 973.607, 51.991783, 3.4127858, 0.18271509, 947.8063, 51.21045, 3.3704734, 0.18242595, 922.39703, 50.426044, 3.3275983, 0.18202724, 897.3806, 49.639202, 3.2842112, 0.18152353, 872.7581, 48.850544, 3.240361, 0.18091933, 848.5303, 48.06067, 3.1960952, 0.18021901, 824.6976, 47.27014, 3.1514597, 0.17942682, 801.2602, 46.479515, 3.1064985, 0.17854694, 778.218, 45.68932, 3.0612543, 0.1775834, 755.5707, 44.900063, 3.0157685, 0.17654017, 733.3177, 44.11223, 2.9700809, 0.17542107, 711.4581, 43.326283, 2.9242294, 0.17422986, 689.991, 42.542675, 2.878251, 0.17297018, 668.91504, 41.76183, 2.8321817, 0.17164555, 648.22864, 40.984158, 2.786055, 0.17025945, 627.93024, 40.21005, 2.7399042, 0.1688152, 608.01794, 39.439877, 2.6937606, 0.16731608, 588.4897, 38.673992, 2.6476548, 0.16576526}};
	localparam real hf[0:1199] = {0.013929818, -9.817731e-06, -1.274517e-05, 1.7709889e-08, 0.013920002, -2.9439356e-05, -1.2708581e-05, 5.3061083e-08, 0.013900385, -4.9019527e-05, -1.2635506e-05, 8.820937e-08, 0.013870994, -6.853073e-05, -1.2526143e-05, 1.2302557e-07, 0.013831871, -8.7945606e-05, -1.2380778e-05, 1.5738583e-07, 0.013783069, -0.000107237, -1.2199782e-05, 1.9117164e-07, 0.013724659, -0.00012637803, -1.1983612e-05, 2.2426991e-07, 0.0136567205, -0.00014534211, -1.1732805e-05, 2.5657306e-07, 0.01357935, -0.0001641031, -1.1447975e-05, 2.87979e-07, 0.013492655, -0.00018263517, -1.112981e-05, 3.1839113e-07, 0.013396757, -0.00020091304, -1.077907e-05, 3.4771847e-07, 0.013291788, -0.00021891196, -1.0396582e-05, 3.7587557e-07, 0.013177896, -0.00023660767, -9.983238e-06, 4.0278252e-07, 0.013055235, -0.00025397656, -9.539991e-06, 4.2836504e-07, 0.012923977, -0.0002709957, -9.067852e-06, 4.525543e-07, 0.012784301, -0.00028764273, -8.567887e-06, 4.75287e-07, 0.0126364, -0.0003038962, -8.04121e-06, 4.965054e-07, 0.012480475, -0.00031973523, -7.488987e-06, 5.16157e-07, 0.012316737, -0.00033513983, -6.9124253e-06, 5.341949e-07, 0.01214541, -0.00035009082, -6.3127727e-06, 5.5057745e-07, 0.011966725, -0.00036456986, -5.6913154e-06, 5.652682e-07, 0.011780922, -0.00037855946, -5.0493727e-06, 5.78236e-07, 0.01158825, -0.0003920431, -4.388294e-06, 5.8945466e-07, 0.011388966, -0.0004050051, -3.709456e-06, 5.9890317e-07, 0.0111833345, -0.00041743074, -3.0142587e-06, 6.0656544e-07, 0.010971626, -0.00042930635, -2.3041223e-06, 6.124301e-07, 0.0107541215, -0.00044061913, -1.580484e-06, 6.1649064e-07, 0.010531103, -0.0004513573, -8.447941e-07, 6.187451e-07, 0.010302862, -0.00046151012, -9.8513596e-08, 6.1919616e-07, 0.0100696925, -0.0004710678, 6.568895e-07, 6.178506e-07, 0.009831894, -0.00048002158, 1.4199431e-06, 6.1471985e-07, 0.009589773, -0.0004883638, 2.1891747e-06, 6.098192e-07, 0.009343633, -0.00049608777, 2.963113e-06, 6.031681e-07, 0.009093788, -0.0005031877, 3.7402924e-06, 5.947897e-07, 0.008840551, -0.0005096591, 4.5192555e-06, 5.847111e-07, 0.008584235, -0.0005154984, 5.2985547e-06, 5.729628e-07, 0.008325159, -0.0005207028, 6.0767566e-06, 5.5957884e-07, 0.008063639, -0.00052527094, 6.8524437e-06, 5.445965e-07, 0.0077999937, -0.0005292021, 7.6242177e-06, 5.2805626e-07, 0.007534542, -0.00053249684, 8.3907e-06, 5.1000154e-07, 0.0072676027, -0.00053515646, 9.150538e-06, 4.904786e-07, 0.0069994912, -0.0005371834, 9.902402e-06, 4.6953633e-07, 0.006730524, -0.00053858105, 1.0644993e-05, 4.4722623e-07, 0.0064610145, -0.0005393537, 1.1377041e-05, 4.2360205e-07, 0.0061912737, -0.0005395065, 1.2097309e-05, 3.9871978e-07, 0.00592161, -0.00053904555, 1.2804592e-05, 3.7263746e-07, 0.005652329, -0.00053797796, 1.34977245e-05, 3.45415e-07, 0.005383732, -0.00053631153, 1.4175575e-05, 3.17114e-07, 0.005116116, -0.00053405494, 1.4837055e-05, 2.877976e-07, 0.004849774, -0.0005312178, 1.5481113e-05, 2.575304e-07, 0.0045849932, -0.00052781036, 1.6106742e-05, 2.263781e-07, 0.0043220567, -0.00052384374, 1.671298e-05, 1.9440763e-07, 0.0040612407, -0.0005193297, 1.7298908e-05, 1.6168676e-07, 0.0038028162, -0.0005142808, 1.7863651e-05, 1.2828403e-07, 0.003547047, -0.0005087103, 1.8406385e-05, 9.426859e-08, 0.0032941906, -0.0005026319, 1.892633e-05, 5.9710075e-08, 0.0030444972, -0.0004960602, 1.9422756e-05, 2.467841e-08, 0.0027982101, -0.00048901024, 1.9894986e-05, -1.07563105e-08, 0.002555564, -0.0004814976, 2.0342386e-05, -4.6523958e-08, 0.002316787, -0.00047353844, 2.0764375e-05, -8.255453e-08, 0.0020820973, -0.00046514938, 2.1160427e-05, -1.1877827e-07, 0.0018517063, -0.0004563475, 2.1530062e-05, -1.5512582e-07, 0.0016258158, -0.00044715032, 2.1872853e-05, -1.9152833e-07, 0.0014046188, -0.00043757574, 2.2188422e-05, -2.279176e-07, 0.0011882999, -0.00042764196, 2.2476446e-05, -2.642262e-07, 0.0009770337, -0.0004173676, 2.2736649e-05, -3.0038763e-07, 0.0007709859, -0.00040677155, 2.2968812e-05, -3.3633629e-07, 0.0005703126, -0.00039587283, 2.317276e-05, -3.720078e-07, 0.0003751603, -0.00038469082, 2.3348373e-05, -4.07339e-07, 0.00018566578, -0.000373245, 2.3495579e-05, -4.4226798e-07, 1.955998e-06, -0.00036155508, 2.3614355e-05, -4.7673433e-07, -0.00017585189, -0.0003496408, 2.3704726e-05, -5.106791e-07, -0.0003476507, -0.00033752198, 2.3766768e-05, -5.4404506e-07, -0.0005133431, -0.0003252186, 2.3800603e-05, -5.7677653e-07, -0.0006728418, -0.00031275052, 2.3806397e-05, -6.0881973e-07, -0.0008260695, -0.00030013768, 2.3784363e-05, -6.4012266e-07, -0.00097295863, -0.0002873999, 2.3734761e-05, -6.7063525e-07, -0.0011134518, -0.00027455695, 2.3657893e-05, -7.0030944e-07, -0.0012475014, -0.00026162853, 2.3554097e-05, -7.2909927e-07, -0.0013750694, -0.00024863417, 2.3423763e-05, -7.5696073e-07, -0.0014961277, -0.00023559315, 2.3267314e-05, -7.8385216e-07, -0.0016106579, -0.00022252469, 2.3085215e-05, -8.0973393e-07, -0.0017186509, -0.00020944767, 2.2877963e-05, -8.345688e-07, -0.0018201072, -0.00019638076, 2.2646096e-05, -8.5832176e-07, -0.0019150365, -0.00018334234, 2.2390188e-05, -8.809601e-07, -0.0020034574, -0.00017035053, 2.211084e-05, -9.0245345e-07, -0.0020853977, -0.00015742303, 2.180869e-05, -9.227738e-07, -0.002160894, -0.00014457724, 2.1484402e-05, -9.4189556e-07, -0.0022299914, -0.00013183017, 2.1138672e-05, -9.597956e-07, -0.0022927434, -0.000119198434, 2.0772222e-05, -9.76453e-07, -0.0023492118, -0.000106698215, 2.0385798e-05, -9.918493e-07, -0.0023994662, -9.434525e-05, 1.9980173e-05, -1.0059688e-06, -0.0024435841, -8.215483e-05, 1.9556135e-05, -1.0187977e-06, -0.0024816506, -7.014176e-05, 1.91145e-05, -1.0303248e-06, -0.0025137577, -5.8320344e-05, 1.8656101e-05, -1.0405414e-06, -0.0025400051, -4.670438e-05, 1.8181787e-05, -1.049441e-06, -0.0025604987, -3.5307137e-05, 1.769242e-05, -1.0570195e-06, -0.0025753507, -2.4141347e-05, 1.718888e-05, -1.0632752e-06, -0.0025846804, -1.3219191e-05, 1.6672058e-05, -1.0682086e-06, -0.0025886125, -2.5522797e-06, 1.6142854e-05, -1.0718223e-06, -0.0025872772, 7.8483445e-06, 1.5602178e-05, -1.0741215e-06, -0.0025808103, 1.7972225e-05, 1.5050946e-05, -1.0751135e-06, -0.0025693527, 2.7809498e-05, 1.4490081e-05, -1.0748072e-06, -0.0025530502, 3.7350892e-05, 1.39205085e-05, -1.0732143e-06, -0.0025320526, 4.658775e-05, 1.3343156e-05, -1.0703483e-06, -0.0025065145, 5.5512013e-05, 1.2758954e-05, -1.0662245e-06, -0.002476594, 6.411625e-05, 1.2168828e-05, -1.0608604e-06, -0.0024424526, 7.2393625e-05, 1.1573705e-05, -1.0542751e-06, -0.0024042558, 8.033794e-05, 1.0974505e-05, -1.04649e-06, -0.0023621712, 8.794359e-05, 1.0372146e-05, -1.0375276e-06, -0.0023163694, 9.520562e-05, 9.767535e-06, -1.0274126e-06, -0.0022670235, 0.000102119666, 9.161573e-06, -1.0161713e-06, -0.0022143084, 0.00010868198, 8.555151e-06, -1.0038314e-06, -0.0021584006, 0.00011488945, 7.949148e-06, -9.904219e-07, -0.0020994786, 0.000120739525, 7.344433e-06, -9.759738e-07, -0.002037721, 0.00012623028, 6.7418578e-06, -9.605187e-07, -0.0019733084, 0.0001313604, 6.1422616e-06, -9.4409035e-07, -0.0019064209, 0.00013612914, 5.546467e-06, -9.26723e-07, -0.0018372395, 0.0001405363, 4.9552796e-06, -9.084522e-07, -0.0017659448, 0.00014458231, 4.3694868e-06, -8.8931466e-07, -0.0016927172, 0.00014826814, 3.789856e-06, -8.693481e-07, -0.0016177364, 0.0001515953, 3.2171347e-06, -8.4859096e-07, -0.0015411814, 0.00015456583, 2.652049e-06, -8.270826e-07, -0.0014632297, 0.00015718232, 2.0953028e-06, -8.0486313e-07, -0.0013840576, 0.00015944787, 1.5475773e-06, -7.819732e-07, -0.0013038396, 0.00016136606, 1.0095295e-06, -7.584542e-07, -0.0012227487, 0.000162941, 4.8179186e-07, -7.343479e-07, -0.0011409551, 0.00016417723, -3.5028133e-08, -7.096966e-07, -0.001058627, 0.00016507978, -5.4034905e-07, -6.8454284e-07, -0.0009759301, 0.0001656541, -1.033616e-06, -6.589295e-07, -0.0008930267, 0.00016590607, -1.5143007e-06, -6.328996e-07, -0.00081007666, 0.00016584201, -1.9819029e-06, -6.0649637e-07, -0.0007272363, 0.00016546859, -2.4359497e-06, -5.79763e-07, -0.00064465846, 0.00016479289, -2.8759966e-06, -5.527427e-07, -0.0005624925, 0.00016382232, -3.3016279e-06, -5.2547847e-07, -0.00048088402, 0.00016256467, -3.7124564e-06, -4.9801326e-07, -0.00039997438, 0.00016102802, -4.1081244e-06, -4.7038975e-07, -0.0003199011, 0.00015922076, -4.4883022e-06, -4.4265033e-07, -0.0002407973, 0.00015715157, -4.8526913e-06, -4.148369e-07, -0.0001627917, 0.00015482941, -5.201021e-06, -3.869911e-07, -8.600852e-05, 0.00015226347, -5.53305e-06, -3.5915386e-07, -1.0567293e-05, 0.00014946317, -5.848568e-06, -3.3136573e-07, 6.3417196e-05, 0.00014643816, -6.1473916e-06, -3.036665e-07, 0.00013583504, 0.00014319825, -6.429367e-06, -2.7609534e-07, 0.0002065813, 0.00013975345, -6.6943717e-06, -2.486907e-07, 0.00027555603, 0.0001361139, -6.9423086e-06, -2.2149014e-07, 0.00034266445, 0.00013228989, -7.17311e-06, -1.945305e-07, 0.0004078169, 0.00012829181, -7.386738e-06, -1.6784766e-07, 0.000470929, 0.00012413017, -7.5831804e-06, -1.4147656e-07, 0.00053192157, 0.00011981552, -7.762452e-06, -1.1545117e-07, 0.0005907208, 0.0001153585, -7.9245965e-06, -8.9804445e-08, 0.00064725813, 0.00011076978, -8.069683e-06, -6.456825e-08, 0.00070147036, 0.00010606005, -8.197805e-06, -3.9773365e-08, 0.00075329974, 0.00010124, -8.309084e-06, -1.5449425e-08, 0.0008026938, 9.632031e-05, -8.403664e-06, 8.375101e-09, 0.00084960525, 9.131164e-05, -8.481714e-06, 3.1672947e-08, 0.0008939923, 8.622457e-05, -8.543426e-06, 5.441807e-08, 0.0009358185, 8.106966e-05, -8.589016e-06, 7.6585685e-08, 0.0009750524, 7.585735e-05, -8.61872e-06, 9.8152285e-08, 0.001011668, 7.0598006e-05, -8.632798e-06, 1.1909564e-07, 0.0010456443, 6.530188e-05, -8.6315285e-06, 1.3939484e-07, 0.0010769655, 5.997908e-05, -8.61521e-06, 1.5903034e-07, 0.0011056205, 5.4639593e-05, -8.584161e-06, 1.7798386e-07, 0.0011316038, 4.9293238e-05, -8.538717e-06, 1.9623855e-07, 0.0011549143, 4.3949673e-05, -8.479233e-06, 2.1377883e-07, 0.0011755556, 3.8618367e-05, -8.406077e-06, 2.3059057e-07, 0.0011935362, 3.33086e-05, -8.3196355e-06, 2.4666096e-07, 0.0012088693, 2.8029439e-05, -8.220309e-06, 2.6197858e-07, 0.0012215723, 2.2789734e-05, -8.108512e-06, 2.7653334e-07, 0.001231667, 1.7598113e-05, -7.98467e-06, 2.903165e-07, 0.0012391797, 1.2462954e-05, -7.849226e-06, 3.0332077e-07, 0.0012441408, 7.3923943e-06, -7.702626e-06, 3.1554012e-07, 0.0012465842, 2.3943069e-06, -7.5453345e-06, 3.2696983e-07, 0.0012465484, -2.5236993e-06, -7.3778197e-06, 3.376066e-07, 0.0012440751, -7.354292e-06, -7.2005605e-06, 3.4744838e-07, 0.0012392098, -1.20904215e-05, -7.0140422e-06, 3.564944e-07, 0.0012320016, -1.6725327e-05, -6.8187587e-06, 3.647452e-07, 0.0012225024, -2.1252545e-05, -6.615207e-06, 3.7220255e-07, 0.001210768, -2.5665911e-05, -6.4038904e-06, 3.7886946e-07, 0.0011968565, -2.9959572e-05, -6.185316e-06, 3.8475014e-07, 0.0011808292, -3.412798e-05, -5.959994e-06, 3.8985e-07, 0.0011627503, -3.816591e-05, -5.728435e-06, 3.9417554e-07, 0.0011426859, -4.206844e-05, -5.491153e-06, 3.977345e-07, 0.0011207052, -4.5830988e-05, -5.248661e-06, 4.0053564e-07, 0.001096879, -4.944929e-05, -5.001473e-06, 4.0258877e-07, 0.0010712806, -5.2919393e-05, -4.750099e-06, 4.0390478e-07, 0.0010439849, -5.6237688e-05, -4.4950493e-06, 4.0449552e-07, 0.0010150687, -5.9400885e-05, -4.2368306e-06, 4.0437385e-07, 0.0009846104, -6.240602e-05, -3.975945e-06, 4.0355349e-07, 0.0009526895, -6.5250446e-05, -3.7128914e-06, 4.020491e-07, 0.0009193871, -6.7931855e-05, -3.4481625e-06, 3.998762e-07, 0.00088478514, -7.044826e-05, -3.1822453e-06, 3.9705108e-07, 0.0008489666, -7.2797986e-05, -2.9156201e-06, 3.9359085e-07, 0.00081201515, -7.4979675e-05, -2.6487603e-06, 3.895133e-07, 0.0007740151, -7.699229e-05, -2.3821303e-06, 3.8483697e-07, 0.0007350512, -7.88351e-05, -2.116187e-06, 3.79581e-07, 0.0006952084, -8.05077e-05, -1.8513771e-06, 3.7376518e-07, 0.00065457186, -8.2009945e-05, -1.5881379e-06, 3.6740985e-07, 0.0006132268, -8.3342034e-05, -1.3268964e-06, 3.6053586e-07, 0.00057125813, -8.450442e-05, -1.0680684e-06, 3.531646e-07, 0.00052875053, -8.549787e-05, -8.1205843e-07, 3.4531783e-07, 0.00048578824, -8.6323416e-05, -5.592591e-07, 3.3701772e-07, 0.00044245488, -8.698236e-05, -3.1005052e-07, 3.2828686e-07, 0.0003988334, -8.747629e-05, -6.48002e-08, 3.1914806e-07, 0.00035500582, -8.780703e-05, 1.7613762e-07, 3.0962445e-07, 0.0003110532, -8.797665e-05, 4.1242225e-07, 2.9973938e-07, 0.0002670556, -8.798751e-05, 6.437268e-07, 2.895164e-07, 0.00022309176, -8.784214e-05, 8.6973876e-07, 2.789792e-07, 0.00017923905, -8.754336e-05, 1.0901599e-06, 2.681515e-07, 0.00013557349, -8.709416e-05, 1.3047066e-06, 2.570572e-07, 9.216944e-05, -8.649776e-05, 1.5131106e-06, 2.4572014e-07, 4.9099683e-05, -8.5757594e-05, 1.7151185e-06, 2.3416418e-07, 6.4352093e-06, -8.487726e-05, 1.9104923e-06, 2.2241308e-07, -3.575484e-05, -8.386055e-05, 2.099009e-06, 2.1049054e-07, -7.740327e-05, -8.2711435e-05, 2.280462e-06, 1.9842012e-07, -0.000118444885, -8.143403e-05, 2.4546596e-06, 1.8622524e-07, -0.00015881662, -8.003263e-05, 2.621426e-06, 1.7392902e-07, -0.00019845758, -7.851165e-05, 2.7806013e-06, 1.6155447e-07, -0.0002373091, -7.687565e-05, 2.9320413e-06, 1.4912422e-07, -0.00027531484, -7.5129305e-05, 3.075617e-06, 1.3666065e-07, -0.0003124208, -7.3277406e-05, 3.211216e-06, 1.2418576e-07, -0.00034857547, -7.132486e-05, 3.3387403e-06, 1.1172124e-07, -0.0003837297, -6.927663e-05, 3.4581083e-06, 9.9288336e-08, -0.000417837, -6.7137815e-05, 3.569253e-06, 8.690786e-08, -0.0004508533, -6.491354e-05, 3.6721235e-06, 7.460021e-08, -0.00048273714, -6.260902e-05, 3.766683e-06, 6.238526e-08, -0.0005134498, -6.02295e-05, 3.85291e-06, 5.0282413e-08, -0.000542955, -5.778029e-05, 3.9307974e-06, 3.8310517e-08, -0.00057121937, -5.5266726e-05, 4.000353e-06, 2.6487884e-08, -0.0005982119, -5.269416e-05, 4.061598e-06, 1.4832247e-08, -0.0006239046, -5.0067967e-05, 4.114567e-06, 3.3607455e-09, -0.0006482718, -4.7393518e-05, 4.1593103e-06, -7.910091e-09, -0.0006712909, -4.467619e-05, 4.1958892e-06, -1.896436e-08, -0.0006929418, -4.1921336e-05, 4.224379e-06, -2.9786808e-08, -0.0007132069, -3.9134295e-05, 4.244867e-06, -4.036283e-08, -0.0007320716, -3.632036e-05, 4.257453e-06, -5.0678512e-08, -0.00074952364, -3.3484805e-05, 4.2622487e-06, -6.07206e-08, -0.0007655536, -3.063284e-05, 4.2593774e-06, -7.047656e-08, -0.0007801546, -2.7769618e-05, 4.248973e-06, -7.993453e-08, -0.0007933222, -2.4900239e-05, 4.2311794e-06, -8.908339e-08, -0.0008050547, -2.202972e-05, 4.2061524e-06, -9.791273e-08, -0.0008153526, -1.9163006e-05, 4.1740564e-06, -1.06412855e-07, -0.0008242191, -1.6304952e-05, 4.135065e-06, -1.145748e-07, -0.00083165977, -1.3460319e-05, 4.0893615e-06, -1.2239033e-07, -0.00083768246, -1.063377e-05, 4.037137e-06, -1.2985194e-07, -0.0008422973, -7.829863e-06, 3.9785905e-06, -1.3695288e-07, -0.0008455168, -5.05304e-06, 3.9139286e-06, -1.4368709e-07, -0.0008473556, -2.3076273e-06, 3.8433654e-06, -1.5004926e-07, -0.0008478304, 4.0217202e-07, 3.7671202e-06, -1.5603482e-07, -0.00084696, 3.0722842e-06, 3.6854199e-06, -1.6163987e-07, -0.00084476534, 5.6987687e-06, 3.5984956e-06, -1.668613e-07, -0.00084126915, 8.277822e-06, 3.5065846e-06, -1.7169664e-07, -0.00083649607, 1.0805785e-05, 3.409928e-06, -1.7614417e-07, -0.00083047245, 1.3279142e-05, 3.3087713e-06, -1.802028e-07, -0.0008232266, 1.5694528e-05, 3.2033633e-06, -1.838722e-07, -0.0008147881, 1.804873e-05, 3.0939566e-06, -1.8715264e-07, -0.00080518855, 2.0338694e-05, 2.9808054e-06, -1.900451e-07, -0.00079446065, 2.256152e-05, 2.8641673e-06, -1.9255116e-07, -0.0007826387, 2.4714473e-05, 2.7443004e-06, -1.9467306e-07, -0.00076975825, 2.6794978e-05, 2.621465e-06, -1.9641367e-07, -0.00075585616, 2.8800627e-05, 2.4959213e-06, -1.9777643e-07, -0.0007409704, 3.0729174e-05, 2.3679306e-06, -1.9876538e-07, -0.00072514015, 3.2578548e-05, 2.2377535e-06, -1.9938514e-07, -0.0007084054, 3.4346835e-05, 2.1056503e-06, -1.9964087e-07, -0.0006908071, 3.6032296e-05, 1.9718802e-06, -1.9953825e-07, -0.0006723872, 3.7633363e-05, 1.8367009e-06, -1.9908352e-07, -0.0006531881, 3.9148632e-05, 1.7003683e-06, -1.9828337e-07, -0.0006332531, 4.057687e-05, 1.5631362e-06, -1.97145e-07, -0.0006126259, 4.1917006e-05, 1.4252553e-06, -1.9567604e-07, -0.0005913509, 4.3168147e-05, 1.2869739e-06, -1.9388457e-07, -0.00056947273, 4.4329554e-05, 1.1485364e-06, -1.917791e-07, -0.00054703635, 4.540066e-05, 1.0101836e-06, -1.8936848e-07, -0.00052408717, 4.638105e-05, 8.721524e-07, -1.8666199e-07, -0.0005006705, 4.727048e-05, 7.3467487e-07, -1.8366924e-07, -0.00047683186, 4.8068865e-05, 5.9797856e-07, -1.8040018e-07, -0.0004526168, 4.877627e-05, 4.6228593e-07, -1.7686502e-07, -0.00042807072, 4.9392907e-05, 3.27814e-07, -1.730743e-07, -0.00040323896, 4.9919156e-05, 1.9477424e-07, -1.690388e-07, -0.00037816656, 5.035553e-05, 6.3372156e-08, -1.6476956e-07, -0.0003528983, 5.070269e-05, -6.61929e-08, -1.6027779e-07, -0.0003274786, 5.0961437e-05, -1.9372797e-07, -1.5557494e-07, -0.00030195143, 5.113271e-05, -3.190467e-07, -1.506726e-07, -0.00027636028, 5.1217583e-05, -4.419696e-07, -1.4558252e-07, -0.00025074807, 5.1217256e-05, -5.623242e-07, -1.4031657e-07, -0.00022515701, 5.1133055e-05, -6.799452e-07, -1.3488673e-07, -0.00019962875, 5.0966424e-05, -7.946746e-07, -1.2930506e-07, -0.00017420408, 5.071893e-05, -9.0636195e-07, -1.2358367e-07, -0.00014892302, 5.0392242e-05, -1.0148646e-06, -1.17734714e-07, -0.00012382474, 4.998815e-05, -1.1200474e-06, -1.11770355e-07, -9.8947465e-05, 4.9508533e-05, -1.2217831e-06, -1.0570276e-07, -7.432846e-05, 4.8955375e-05, -1.3199527e-06, -9.954407e-08, -5.0004e-05, 4.833075e-05, -1.4144447e-06, -9.330637e-08, -2.600927e-05, 4.7636815e-05, -1.5051561e-06, -8.7001695e-08, -2.3783643e-06, 4.6875823e-05, -1.5919919e-06, -8.064199e-08, 2.0855761e-05, 4.6050092e-05, -1.6748651e-06, -7.423908e-08, 4.3661334e-05, 4.5162018e-05, -1.7536969e-06, -6.780471e-08, 6.600779e-05, 4.421406e-05, -1.8284169e-06, -6.135044e-08, 8.786583e-05, 4.3208744e-05, -1.8989624e-06, -5.4887696e-08, 0.00010920741, 4.2148644e-05, -1.9652794e-06, -4.8427726e-08, 0.00013000578, 4.1036394e-05, -2.0273214e-06, -4.1981586e-08};
	localparam real hb[0:1199] = {0.013929818, 9.817731e-06, -1.274517e-05, -1.7709889e-08, 0.013920002, 2.9439356e-05, -1.2708581e-05, -5.3061083e-08, 0.013900385, 4.9019527e-05, -1.2635506e-05, -8.820937e-08, 0.013870994, 6.853073e-05, -1.2526143e-05, -1.2302557e-07, 0.013831871, 8.7945606e-05, -1.2380778e-05, -1.5738583e-07, 0.013783069, 0.000107237, -1.2199782e-05, -1.9117164e-07, 0.013724659, 0.00012637803, -1.1983612e-05, -2.2426991e-07, 0.0136567205, 0.00014534211, -1.1732805e-05, -2.5657306e-07, 0.01357935, 0.0001641031, -1.1447975e-05, -2.87979e-07, 0.013492655, 0.00018263517, -1.112981e-05, -3.1839113e-07, 0.013396757, 0.00020091304, -1.077907e-05, -3.4771847e-07, 0.013291788, 0.00021891196, -1.0396582e-05, -3.7587557e-07, 0.013177896, 0.00023660767, -9.983238e-06, -4.0278252e-07, 0.013055235, 0.00025397656, -9.539991e-06, -4.2836504e-07, 0.012923977, 0.0002709957, -9.067852e-06, -4.525543e-07, 0.012784301, 0.00028764273, -8.567887e-06, -4.75287e-07, 0.0126364, 0.0003038962, -8.04121e-06, -4.965054e-07, 0.012480475, 0.00031973523, -7.488987e-06, -5.16157e-07, 0.012316737, 0.00033513983, -6.9124253e-06, -5.341949e-07, 0.01214541, 0.00035009082, -6.3127727e-06, -5.5057745e-07, 0.011966725, 0.00036456986, -5.6913154e-06, -5.652682e-07, 0.011780922, 0.00037855946, -5.0493727e-06, -5.78236e-07, 0.01158825, 0.0003920431, -4.388294e-06, -5.8945466e-07, 0.011388966, 0.0004050051, -3.709456e-06, -5.9890317e-07, 0.0111833345, 0.00041743074, -3.0142587e-06, -6.0656544e-07, 0.010971626, 0.00042930635, -2.3041223e-06, -6.124301e-07, 0.0107541215, 0.00044061913, -1.580484e-06, -6.1649064e-07, 0.010531103, 0.0004513573, -8.447941e-07, -6.187451e-07, 0.010302862, 0.00046151012, -9.8513596e-08, -6.1919616e-07, 0.0100696925, 0.0004710678, 6.568895e-07, -6.178506e-07, 0.009831894, 0.00048002158, 1.4199431e-06, -6.1471985e-07, 0.009589773, 0.0004883638, 2.1891747e-06, -6.098192e-07, 0.009343633, 0.00049608777, 2.963113e-06, -6.031681e-07, 0.009093788, 0.0005031877, 3.7402924e-06, -5.947897e-07, 0.008840551, 0.0005096591, 4.5192555e-06, -5.847111e-07, 0.008584235, 0.0005154984, 5.2985547e-06, -5.729628e-07, 0.008325159, 0.0005207028, 6.0767566e-06, -5.5957884e-07, 0.008063639, 0.00052527094, 6.8524437e-06, -5.445965e-07, 0.0077999937, 0.0005292021, 7.6242177e-06, -5.2805626e-07, 0.007534542, 0.00053249684, 8.3907e-06, -5.1000154e-07, 0.0072676027, 0.00053515646, 9.150538e-06, -4.904786e-07, 0.0069994912, 0.0005371834, 9.902402e-06, -4.6953633e-07, 0.006730524, 0.00053858105, 1.0644993e-05, -4.4722623e-07, 0.0064610145, 0.0005393537, 1.1377041e-05, -4.2360205e-07, 0.0061912737, 0.0005395065, 1.2097309e-05, -3.9871978e-07, 0.00592161, 0.00053904555, 1.2804592e-05, -3.7263746e-07, 0.005652329, 0.00053797796, 1.34977245e-05, -3.45415e-07, 0.005383732, 0.00053631153, 1.4175575e-05, -3.17114e-07, 0.005116116, 0.00053405494, 1.4837055e-05, -2.877976e-07, 0.004849774, 0.0005312178, 1.5481113e-05, -2.575304e-07, 0.0045849932, 0.00052781036, 1.6106742e-05, -2.263781e-07, 0.0043220567, 0.00052384374, 1.671298e-05, -1.9440763e-07, 0.0040612407, 0.0005193297, 1.7298908e-05, -1.6168676e-07, 0.0038028162, 0.0005142808, 1.7863651e-05, -1.2828403e-07, 0.003547047, 0.0005087103, 1.8406385e-05, -9.426859e-08, 0.0032941906, 0.0005026319, 1.892633e-05, -5.9710075e-08, 0.0030444972, 0.0004960602, 1.9422756e-05, -2.467841e-08, 0.0027982101, 0.00048901024, 1.9894986e-05, 1.07563105e-08, 0.002555564, 0.0004814976, 2.0342386e-05, 4.6523958e-08, 0.002316787, 0.00047353844, 2.0764375e-05, 8.255453e-08, 0.0020820973, 0.00046514938, 2.1160427e-05, 1.1877827e-07, 0.0018517063, 0.0004563475, 2.1530062e-05, 1.5512582e-07, 0.0016258158, 0.00044715032, 2.1872853e-05, 1.9152833e-07, 0.0014046188, 0.00043757574, 2.2188422e-05, 2.279176e-07, 0.0011882999, 0.00042764196, 2.2476446e-05, 2.642262e-07, 0.0009770337, 0.0004173676, 2.2736649e-05, 3.0038763e-07, 0.0007709859, 0.00040677155, 2.2968812e-05, 3.3633629e-07, 0.0005703126, 0.00039587283, 2.317276e-05, 3.720078e-07, 0.0003751603, 0.00038469082, 2.3348373e-05, 4.07339e-07, 0.00018566578, 0.000373245, 2.3495579e-05, 4.4226798e-07, 1.955998e-06, 0.00036155508, 2.3614355e-05, 4.7673433e-07, -0.00017585189, 0.0003496408, 2.3704726e-05, 5.106791e-07, -0.0003476507, 0.00033752198, 2.3766768e-05, 5.4404506e-07, -0.0005133431, 0.0003252186, 2.3800603e-05, 5.7677653e-07, -0.0006728418, 0.00031275052, 2.3806397e-05, 6.0881973e-07, -0.0008260695, 0.00030013768, 2.3784363e-05, 6.4012266e-07, -0.00097295863, 0.0002873999, 2.3734761e-05, 6.7063525e-07, -0.0011134518, 0.00027455695, 2.3657893e-05, 7.0030944e-07, -0.0012475014, 0.00026162853, 2.3554097e-05, 7.2909927e-07, -0.0013750694, 0.00024863417, 2.3423763e-05, 7.5696073e-07, -0.0014961277, 0.00023559315, 2.3267314e-05, 7.8385216e-07, -0.0016106579, 0.00022252469, 2.3085215e-05, 8.0973393e-07, -0.0017186509, 0.00020944767, 2.2877963e-05, 8.345688e-07, -0.0018201072, 0.00019638076, 2.2646096e-05, 8.5832176e-07, -0.0019150365, 0.00018334234, 2.2390188e-05, 8.809601e-07, -0.0020034574, 0.00017035053, 2.211084e-05, 9.0245345e-07, -0.0020853977, 0.00015742303, 2.180869e-05, 9.227738e-07, -0.002160894, 0.00014457724, 2.1484402e-05, 9.4189556e-07, -0.0022299914, 0.00013183017, 2.1138672e-05, 9.597956e-07, -0.0022927434, 0.000119198434, 2.0772222e-05, 9.76453e-07, -0.0023492118, 0.000106698215, 2.0385798e-05, 9.918493e-07, -0.0023994662, 9.434525e-05, 1.9980173e-05, 1.0059688e-06, -0.0024435841, 8.215483e-05, 1.9556135e-05, 1.0187977e-06, -0.0024816506, 7.014176e-05, 1.91145e-05, 1.0303248e-06, -0.0025137577, 5.8320344e-05, 1.8656101e-05, 1.0405414e-06, -0.0025400051, 4.670438e-05, 1.8181787e-05, 1.049441e-06, -0.0025604987, 3.5307137e-05, 1.769242e-05, 1.0570195e-06, -0.0025753507, 2.4141347e-05, 1.718888e-05, 1.0632752e-06, -0.0025846804, 1.3219191e-05, 1.6672058e-05, 1.0682086e-06, -0.0025886125, 2.5522797e-06, 1.6142854e-05, 1.0718223e-06, -0.0025872772, -7.8483445e-06, 1.5602178e-05, 1.0741215e-06, -0.0025808103, -1.7972225e-05, 1.5050946e-05, 1.0751135e-06, -0.0025693527, -2.7809498e-05, 1.4490081e-05, 1.0748072e-06, -0.0025530502, -3.7350892e-05, 1.39205085e-05, 1.0732143e-06, -0.0025320526, -4.658775e-05, 1.3343156e-05, 1.0703483e-06, -0.0025065145, -5.5512013e-05, 1.2758954e-05, 1.0662245e-06, -0.002476594, -6.411625e-05, 1.2168828e-05, 1.0608604e-06, -0.0024424526, -7.2393625e-05, 1.1573705e-05, 1.0542751e-06, -0.0024042558, -8.033794e-05, 1.0974505e-05, 1.04649e-06, -0.0023621712, -8.794359e-05, 1.0372146e-05, 1.0375276e-06, -0.0023163694, -9.520562e-05, 9.767535e-06, 1.0274126e-06, -0.0022670235, -0.000102119666, 9.161573e-06, 1.0161713e-06, -0.0022143084, -0.00010868198, 8.555151e-06, 1.0038314e-06, -0.0021584006, -0.00011488945, 7.949148e-06, 9.904219e-07, -0.0020994786, -0.000120739525, 7.344433e-06, 9.759738e-07, -0.002037721, -0.00012623028, 6.7418578e-06, 9.605187e-07, -0.0019733084, -0.0001313604, 6.1422616e-06, 9.4409035e-07, -0.0019064209, -0.00013612914, 5.546467e-06, 9.26723e-07, -0.0018372395, -0.0001405363, 4.9552796e-06, 9.084522e-07, -0.0017659448, -0.00014458231, 4.3694868e-06, 8.8931466e-07, -0.0016927172, -0.00014826814, 3.789856e-06, 8.693481e-07, -0.0016177364, -0.0001515953, 3.2171347e-06, 8.4859096e-07, -0.0015411814, -0.00015456583, 2.652049e-06, 8.270826e-07, -0.0014632297, -0.00015718232, 2.0953028e-06, 8.0486313e-07, -0.0013840576, -0.00015944787, 1.5475773e-06, 7.819732e-07, -0.0013038396, -0.00016136606, 1.0095295e-06, 7.584542e-07, -0.0012227487, -0.000162941, 4.8179186e-07, 7.343479e-07, -0.0011409551, -0.00016417723, -3.5028133e-08, 7.096966e-07, -0.001058627, -0.00016507978, -5.4034905e-07, 6.8454284e-07, -0.0009759301, -0.0001656541, -1.033616e-06, 6.589295e-07, -0.0008930267, -0.00016590607, -1.5143007e-06, 6.328996e-07, -0.00081007666, -0.00016584201, -1.9819029e-06, 6.0649637e-07, -0.0007272363, -0.00016546859, -2.4359497e-06, 5.79763e-07, -0.00064465846, -0.00016479289, -2.8759966e-06, 5.527427e-07, -0.0005624925, -0.00016382232, -3.3016279e-06, 5.2547847e-07, -0.00048088402, -0.00016256467, -3.7124564e-06, 4.9801326e-07, -0.00039997438, -0.00016102802, -4.1081244e-06, 4.7038975e-07, -0.0003199011, -0.00015922076, -4.4883022e-06, 4.4265033e-07, -0.0002407973, -0.00015715157, -4.8526913e-06, 4.148369e-07, -0.0001627917, -0.00015482941, -5.201021e-06, 3.869911e-07, -8.600852e-05, -0.00015226347, -5.53305e-06, 3.5915386e-07, -1.0567293e-05, -0.00014946317, -5.848568e-06, 3.3136573e-07, 6.3417196e-05, -0.00014643816, -6.1473916e-06, 3.036665e-07, 0.00013583504, -0.00014319825, -6.429367e-06, 2.7609534e-07, 0.0002065813, -0.00013975345, -6.6943717e-06, 2.486907e-07, 0.00027555603, -0.0001361139, -6.9423086e-06, 2.2149014e-07, 0.00034266445, -0.00013228989, -7.17311e-06, 1.945305e-07, 0.0004078169, -0.00012829181, -7.386738e-06, 1.6784766e-07, 0.000470929, -0.00012413017, -7.5831804e-06, 1.4147656e-07, 0.00053192157, -0.00011981552, -7.762452e-06, 1.1545117e-07, 0.0005907208, -0.0001153585, -7.9245965e-06, 8.9804445e-08, 0.00064725813, -0.00011076978, -8.069683e-06, 6.456825e-08, 0.00070147036, -0.00010606005, -8.197805e-06, 3.9773365e-08, 0.00075329974, -0.00010124, -8.309084e-06, 1.5449425e-08, 0.0008026938, -9.632031e-05, -8.403664e-06, -8.375101e-09, 0.00084960525, -9.131164e-05, -8.481714e-06, -3.1672947e-08, 0.0008939923, -8.622457e-05, -8.543426e-06, -5.441807e-08, 0.0009358185, -8.106966e-05, -8.589016e-06, -7.6585685e-08, 0.0009750524, -7.585735e-05, -8.61872e-06, -9.8152285e-08, 0.001011668, -7.0598006e-05, -8.632798e-06, -1.1909564e-07, 0.0010456443, -6.530188e-05, -8.6315285e-06, -1.3939484e-07, 0.0010769655, -5.997908e-05, -8.61521e-06, -1.5903034e-07, 0.0011056205, -5.4639593e-05, -8.584161e-06, -1.7798386e-07, 0.0011316038, -4.9293238e-05, -8.538717e-06, -1.9623855e-07, 0.0011549143, -4.3949673e-05, -8.479233e-06, -2.1377883e-07, 0.0011755556, -3.8618367e-05, -8.406077e-06, -2.3059057e-07, 0.0011935362, -3.33086e-05, -8.3196355e-06, -2.4666096e-07, 0.0012088693, -2.8029439e-05, -8.220309e-06, -2.6197858e-07, 0.0012215723, -2.2789734e-05, -8.108512e-06, -2.7653334e-07, 0.001231667, -1.7598113e-05, -7.98467e-06, -2.903165e-07, 0.0012391797, -1.2462954e-05, -7.849226e-06, -3.0332077e-07, 0.0012441408, -7.3923943e-06, -7.702626e-06, -3.1554012e-07, 0.0012465842, -2.3943069e-06, -7.5453345e-06, -3.2696983e-07, 0.0012465484, 2.5236993e-06, -7.3778197e-06, -3.376066e-07, 0.0012440751, 7.354292e-06, -7.2005605e-06, -3.4744838e-07, 0.0012392098, 1.20904215e-05, -7.0140422e-06, -3.564944e-07, 0.0012320016, 1.6725327e-05, -6.8187587e-06, -3.647452e-07, 0.0012225024, 2.1252545e-05, -6.615207e-06, -3.7220255e-07, 0.001210768, 2.5665911e-05, -6.4038904e-06, -3.7886946e-07, 0.0011968565, 2.9959572e-05, -6.185316e-06, -3.8475014e-07, 0.0011808292, 3.412798e-05, -5.959994e-06, -3.8985e-07, 0.0011627503, 3.816591e-05, -5.728435e-06, -3.9417554e-07, 0.0011426859, 4.206844e-05, -5.491153e-06, -3.977345e-07, 0.0011207052, 4.5830988e-05, -5.248661e-06, -4.0053564e-07, 0.001096879, 4.944929e-05, -5.001473e-06, -4.0258877e-07, 0.0010712806, 5.2919393e-05, -4.750099e-06, -4.0390478e-07, 0.0010439849, 5.6237688e-05, -4.4950493e-06, -4.0449552e-07, 0.0010150687, 5.9400885e-05, -4.2368306e-06, -4.0437385e-07, 0.0009846104, 6.240602e-05, -3.975945e-06, -4.0355349e-07, 0.0009526895, 6.5250446e-05, -3.7128914e-06, -4.020491e-07, 0.0009193871, 6.7931855e-05, -3.4481625e-06, -3.998762e-07, 0.00088478514, 7.044826e-05, -3.1822453e-06, -3.9705108e-07, 0.0008489666, 7.2797986e-05, -2.9156201e-06, -3.9359085e-07, 0.00081201515, 7.4979675e-05, -2.6487603e-06, -3.895133e-07, 0.0007740151, 7.699229e-05, -2.3821303e-06, -3.8483697e-07, 0.0007350512, 7.88351e-05, -2.116187e-06, -3.79581e-07, 0.0006952084, 8.05077e-05, -1.8513771e-06, -3.7376518e-07, 0.00065457186, 8.2009945e-05, -1.5881379e-06, -3.6740985e-07, 0.0006132268, 8.3342034e-05, -1.3268964e-06, -3.6053586e-07, 0.00057125813, 8.450442e-05, -1.0680684e-06, -3.531646e-07, 0.00052875053, 8.549787e-05, -8.1205843e-07, -3.4531783e-07, 0.00048578824, 8.6323416e-05, -5.592591e-07, -3.3701772e-07, 0.00044245488, 8.698236e-05, -3.1005052e-07, -3.2828686e-07, 0.0003988334, 8.747629e-05, -6.48002e-08, -3.1914806e-07, 0.00035500582, 8.780703e-05, 1.7613762e-07, -3.0962445e-07, 0.0003110532, 8.797665e-05, 4.1242225e-07, -2.9973938e-07, 0.0002670556, 8.798751e-05, 6.437268e-07, -2.895164e-07, 0.00022309176, 8.784214e-05, 8.6973876e-07, -2.789792e-07, 0.00017923905, 8.754336e-05, 1.0901599e-06, -2.681515e-07, 0.00013557349, 8.709416e-05, 1.3047066e-06, -2.570572e-07, 9.216944e-05, 8.649776e-05, 1.5131106e-06, -2.4572014e-07, 4.9099683e-05, 8.5757594e-05, 1.7151185e-06, -2.3416418e-07, 6.4352093e-06, 8.487726e-05, 1.9104923e-06, -2.2241308e-07, -3.575484e-05, 8.386055e-05, 2.099009e-06, -2.1049054e-07, -7.740327e-05, 8.2711435e-05, 2.280462e-06, -1.9842012e-07, -0.000118444885, 8.143403e-05, 2.4546596e-06, -1.8622524e-07, -0.00015881662, 8.003263e-05, 2.621426e-06, -1.7392902e-07, -0.00019845758, 7.851165e-05, 2.7806013e-06, -1.6155447e-07, -0.0002373091, 7.687565e-05, 2.9320413e-06, -1.4912422e-07, -0.00027531484, 7.5129305e-05, 3.075617e-06, -1.3666065e-07, -0.0003124208, 7.3277406e-05, 3.211216e-06, -1.2418576e-07, -0.00034857547, 7.132486e-05, 3.3387403e-06, -1.1172124e-07, -0.0003837297, 6.927663e-05, 3.4581083e-06, -9.9288336e-08, -0.000417837, 6.7137815e-05, 3.569253e-06, -8.690786e-08, -0.0004508533, 6.491354e-05, 3.6721235e-06, -7.460021e-08, -0.00048273714, 6.260902e-05, 3.766683e-06, -6.238526e-08, -0.0005134498, 6.02295e-05, 3.85291e-06, -5.0282413e-08, -0.000542955, 5.778029e-05, 3.9307974e-06, -3.8310517e-08, -0.00057121937, 5.5266726e-05, 4.000353e-06, -2.6487884e-08, -0.0005982119, 5.269416e-05, 4.061598e-06, -1.4832247e-08, -0.0006239046, 5.0067967e-05, 4.114567e-06, -3.3607455e-09, -0.0006482718, 4.7393518e-05, 4.1593103e-06, 7.910091e-09, -0.0006712909, 4.467619e-05, 4.1958892e-06, 1.896436e-08, -0.0006929418, 4.1921336e-05, 4.224379e-06, 2.9786808e-08, -0.0007132069, 3.9134295e-05, 4.244867e-06, 4.036283e-08, -0.0007320716, 3.632036e-05, 4.257453e-06, 5.0678512e-08, -0.00074952364, 3.3484805e-05, 4.2622487e-06, 6.07206e-08, -0.0007655536, 3.063284e-05, 4.2593774e-06, 7.047656e-08, -0.0007801546, 2.7769618e-05, 4.248973e-06, 7.993453e-08, -0.0007933222, 2.4900239e-05, 4.2311794e-06, 8.908339e-08, -0.0008050547, 2.202972e-05, 4.2061524e-06, 9.791273e-08, -0.0008153526, 1.9163006e-05, 4.1740564e-06, 1.06412855e-07, -0.0008242191, 1.6304952e-05, 4.135065e-06, 1.145748e-07, -0.00083165977, 1.3460319e-05, 4.0893615e-06, 1.2239033e-07, -0.00083768246, 1.063377e-05, 4.037137e-06, 1.2985194e-07, -0.0008422973, 7.829863e-06, 3.9785905e-06, 1.3695288e-07, -0.0008455168, 5.05304e-06, 3.9139286e-06, 1.4368709e-07, -0.0008473556, 2.3076273e-06, 3.8433654e-06, 1.5004926e-07, -0.0008478304, -4.0217202e-07, 3.7671202e-06, 1.5603482e-07, -0.00084696, -3.0722842e-06, 3.6854199e-06, 1.6163987e-07, -0.00084476534, -5.6987687e-06, 3.5984956e-06, 1.668613e-07, -0.00084126915, -8.277822e-06, 3.5065846e-06, 1.7169664e-07, -0.00083649607, -1.0805785e-05, 3.409928e-06, 1.7614417e-07, -0.00083047245, -1.3279142e-05, 3.3087713e-06, 1.802028e-07, -0.0008232266, -1.5694528e-05, 3.2033633e-06, 1.838722e-07, -0.0008147881, -1.804873e-05, 3.0939566e-06, 1.8715264e-07, -0.00080518855, -2.0338694e-05, 2.9808054e-06, 1.900451e-07, -0.00079446065, -2.256152e-05, 2.8641673e-06, 1.9255116e-07, -0.0007826387, -2.4714473e-05, 2.7443004e-06, 1.9467306e-07, -0.00076975825, -2.6794978e-05, 2.621465e-06, 1.9641367e-07, -0.00075585616, -2.8800627e-05, 2.4959213e-06, 1.9777643e-07, -0.0007409704, -3.0729174e-05, 2.3679306e-06, 1.9876538e-07, -0.00072514015, -3.2578548e-05, 2.2377535e-06, 1.9938514e-07, -0.0007084054, -3.4346835e-05, 2.1056503e-06, 1.9964087e-07, -0.0006908071, -3.6032296e-05, 1.9718802e-06, 1.9953825e-07, -0.0006723872, -3.7633363e-05, 1.8367009e-06, 1.9908352e-07, -0.0006531881, -3.9148632e-05, 1.7003683e-06, 1.9828337e-07, -0.0006332531, -4.057687e-05, 1.5631362e-06, 1.97145e-07, -0.0006126259, -4.1917006e-05, 1.4252553e-06, 1.9567604e-07, -0.0005913509, -4.3168147e-05, 1.2869739e-06, 1.9388457e-07, -0.00056947273, -4.4329554e-05, 1.1485364e-06, 1.917791e-07, -0.00054703635, -4.540066e-05, 1.0101836e-06, 1.8936848e-07, -0.00052408717, -4.638105e-05, 8.721524e-07, 1.8666199e-07, -0.0005006705, -4.727048e-05, 7.3467487e-07, 1.8366924e-07, -0.00047683186, -4.8068865e-05, 5.9797856e-07, 1.8040018e-07, -0.0004526168, -4.877627e-05, 4.6228593e-07, 1.7686502e-07, -0.00042807072, -4.9392907e-05, 3.27814e-07, 1.730743e-07, -0.00040323896, -4.9919156e-05, 1.9477424e-07, 1.690388e-07, -0.00037816656, -5.035553e-05, 6.3372156e-08, 1.6476956e-07, -0.0003528983, -5.070269e-05, -6.61929e-08, 1.6027779e-07, -0.0003274786, -5.0961437e-05, -1.9372797e-07, 1.5557494e-07, -0.00030195143, -5.113271e-05, -3.190467e-07, 1.506726e-07, -0.00027636028, -5.1217583e-05, -4.419696e-07, 1.4558252e-07, -0.00025074807, -5.1217256e-05, -5.623242e-07, 1.4031657e-07, -0.00022515701, -5.1133055e-05, -6.799452e-07, 1.3488673e-07, -0.00019962875, -5.0966424e-05, -7.946746e-07, 1.2930506e-07, -0.00017420408, -5.071893e-05, -9.0636195e-07, 1.2358367e-07, -0.00014892302, -5.0392242e-05, -1.0148646e-06, 1.17734714e-07, -0.00012382474, -4.998815e-05, -1.1200474e-06, 1.11770355e-07, -9.8947465e-05, -4.9508533e-05, -1.2217831e-06, 1.0570276e-07, -7.432846e-05, -4.8955375e-05, -1.3199527e-06, 9.954407e-08, -5.0004e-05, -4.833075e-05, -1.4144447e-06, 9.330637e-08, -2.600927e-05, -4.7636815e-05, -1.5051561e-06, 8.7001695e-08, -2.3783643e-06, -4.6875823e-05, -1.5919919e-06, 8.064199e-08, 2.0855761e-05, -4.6050092e-05, -1.6748651e-06, 7.423908e-08, 4.3661334e-05, -4.5162018e-05, -1.7536969e-06, 6.780471e-08, 6.600779e-05, -4.421406e-05, -1.8284169e-06, 6.135044e-08, 8.786583e-05, -4.3208744e-05, -1.8989624e-06, 5.4887696e-08, 0.00010920741, -4.2148644e-05, -1.9652794e-06, 4.8427726e-08, 0.00013000578, -4.1036394e-05, -2.0273214e-06, 4.1981586e-08};
endpackage
`endif
