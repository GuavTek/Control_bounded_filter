`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam N = 4;
	localparam COEFF_BIAS = 48;
	localparam logic signed[63:0] Lfr[0:3] = {64'd277489893271481, 64'd277489893271481, 64'd275315491622285, 64'd275315491622285};
	localparam logic signed[63:0] Lfi[0:3] = {64'd30020001337947, - 64'd30020001337947, 64'd11558098293529, - 64'd11558098293529};
	localparam logic signed[63:0] Lbr[0:3] = {64'd277489893271481, 64'd277489893271481, 64'd275315491622285, 64'd275315491622285};
	localparam logic signed[63:0] Lbi[0:3] = {64'd30020001337947, - 64'd30020001337947, 64'd11558098293529, - 64'd11558098293529};
	localparam logic signed[63:0] Wfr[0:3] = {64'd24193209882, 64'd24193209882, - 64'd7887428590, - 64'd7887428590};
	localparam logic signed[63:0] Wfi[0:3] = {64'd29297075841, - 64'd29297075841, - 64'd33126712469, 64'd33126712469};
	localparam logic signed[63:0] Wbr[0:3] = {- 64'd24193209882, - 64'd24193209882, 64'd7887428590, 64'd7887428590};
	localparam logic signed[63:0] Wbi[0:3] = {- 64'd29297075841, 64'd29297075841, 64'd33126712469, - 64'd33126712469};
	localparam logic signed[63:0] Ffr[0:3][0:79] = '{
		'{64'd2678910912348682, 64'd1633669149297615, - 64'd134405106412023, - 64'd14489081406757, 64'd3471761733289509, 64'd1534935316807140, - 64'd154547576200402, - 64'd12167341321049, 64'd4211153497515380, 64'd1420087166233641, - 64'd172563932222687, - 64'd9743629047954, 64'd4889422534499934, 64'd1290723849399400, - 64'd188281223922595, - 64'd7247706595933, 64'd5499740975037776, 64'd1148585763351890, - 64'd201556008143343, - 64'd4709673588602, 64'd6036181793402482, 64'd995532040410431, - 64'd212275515540637, - 64'd2159613203878, 64'd6493772333226378, 64'd833517040657504, - 64'd220358442413966, 64'd372755769329, 64'd6868535890318197, 64'd664566135678268, - 64'd225755365061278, 64'd2858416831816, 64'd7157521071022570, 64'd490751075721102, - 64'd228448778179966, 64'd5269379888993, 64'd7358818790936519, 64'd314165232382821, - 64'd228452763163329, 64'd7578988059119, 64'd7471566924126414, 64'd136899005473061, - 64'd225812296327788, 64'd9762203913194, 64'd7495942755766966, - 64'd38984324020268, - 64'd220602211106000, 64'd11795872177577, 64'd7433143529741519, - 64'd211472022825834, - 64'd212925832011491, 64'd13658956252499, 64'd7285355515665612, - 64'd378624356972050, - 64'd202913301681643, 64'd15332746247078, 64'd7055712145579892, - 64'd538595822537850, - 64'd190719625501872, 64'd16801036599608, 64'd6748241887867779, - 64'd689654930258371, - 64'd176522461172683, 64'd18050271736293, 64'd6367806633571694, - 64'd830202339184127, - 64'd160519683075600, 64'd19069658617453, 64'd5920031467125635, - 64'd958787157130758, - 64'd142926753400873, 64'd19851245422781, 64'd5411226778650929, - 64'd1074121249927379, - 64'd123973933701595, 64'd20389966031699, 64'd4848303747586724, - 64'd1175091427164946, - 64'd103903371822373, 64'd20683650356549},
		'{64'd2678910912348222, 64'd1633669149297648, - 64'd134405106412032, - 64'd14489081406755, 64'd3471761733289070, 64'd1534935316807172, - 64'd154547576200411, - 64'd12167341321048, 64'd4211153497514966, 64'd1420087166233671, - 64'd172563932222695, - 64'd9743629047952, 64'd4889422534499551, 64'd1290723849399429, - 64'd188281223922603, - 64'd7247706595932, 64'd5499740975037427, 64'd1148585763351916, - 64'd201556008143349, - 64'd4709673588600, 64'd6036181793402171, 64'd995532040410455, - 64'd212275515540643, - 64'd2159613203877, 64'd6493772333226108, 64'd833517040657526, - 64'd220358442413972, 64'd372755769330, 64'd6868535890317968, 64'd664566135678286, - 64'd225755365061283, 64'd2858416831817, 64'd7157521071022387, 64'd490751075721118, - 64'd228448778179969, 64'd5269379888994, 64'd7358818790936382, 64'd314165232382833, - 64'd228452763163332, 64'd7578988059119, 64'd7471566924126326, 64'd136899005473070, - 64'd225812296327790, 64'd9762203913194, 64'd7495942755766923, - 64'd38984324020262, - 64'd220602211106001, 64'd11795872177577, 64'd7433143529741523, - 64'd211472022825831, - 64'd212925832011491, 64'd13658956252499, 64'd7285355515665663, - 64'd378624356972050, - 64'd202913301681642, 64'd15332746247078, 64'd7055712145579987, - 64'd538595822537854, - 64'd190719625501870, 64'd16801036599608, 64'd6748241887867917, - 64'd689654930258378, - 64'd176522461172680, 64'd18050271736292, 64'd6367806633571872, - 64'd830202339184137, - 64'd160519683075597, 64'd19069658617452, 64'd5920031467125852, - 64'd958787157130771, - 64'd142926753400869, 64'd19851245422781, 64'd5411226778651180, - 64'd1074121249927394, - 64'd123973933701590, 64'd20389966031698, 64'd4848303747587006, - 64'd1175091427164964, - 64'd103903371822367, 64'd20683650356548},
		'{- 64'd2621464726625032, - 64'd1601298142322358, 64'd114277463862052, - 64'd54557765512014, - 64'd3402192470904109, - 64'd1521613693668172, 64'd101035526953527, - 64'd52555428834631, - 64'd4143075592769200, - 64'd1441949887694716, 64'd88125723066021, - 64'd50522608463608, - 64'd4844167648167600, - 64'd1362478337710847, 64'd75562184921028, - 64'd48464973598293, - 64'd5505606112696863, - 64'd1283363101544773, 64'd63357707642890, - 64'd46388011318305, - 64'd6127608592847788, - 64'd1204760640672868, 64'd51523776702445, - 64'd44297022280332, - 64'd6710469021379336, - 64'd1126819797494854, 64'd40070597533593, - 64'd42197116997554, - 64'd7254553845722606, - 64'd1049681790049648, 64'd29007126689070, - 64'd40093212685504, - 64'd7760298217955961, - 64'd973480223457764, 64'd18341104403946, - 64'd37990030657633, - 64'd8228202194534652, - 64'd898341117369665, 64'd8079088437780, - 64'd35892094253348, - 64'd8658826953596720, - 64'd824382948694780, - 64'd1773510931025, - 64'd33803727280864, - 64'd9052791037303526, - 64'd751716708882984, - 64'd11212394882364, - 64'd31729052956814, - 64'd9410766626308762, - 64'd680445975029133, - 64'd20234339123843, - 64'd29671993324251, - 64'd9733475853085184, - 64'd610666994071677, - 64'd28837156170190, - 64'd27636269130411, - 64'd10021687160474126, - 64'd542468779358319, - 64'd37019656947170, - 64'd25625400145358, - 64'd10276211711460314, - 64'd475933218855185, - 64'd44781611831263, - 64'd23642705902492, - 64'd10497899855813746, - 64'd411135194280852, - 64'd52123711232903, - 64'd21691306841762, - 64'd10687637658882664, - 64'd348142710452834, - 64'd59047525827614, - 64'd19774125836360, - 64'd10846343497467206, - 64'd287017034141629, - 64'd65555466535792, - 64'd17893890083631, - 64'd10974964727353150, - 64'd227812841736200, - 64'd71650744348225, - 64'd16053133340965},
		'{- 64'd2621464726623828, - 64'd1601298142322414, 64'd114277463862073, - 64'd54557765512018, - 64'd3402192470902937, - 64'd1521613693668227, 64'd101035526953548, - 64'd52555428834635, - 64'd4143075592768060, - 64'd1441949887694769, 64'd88125723066041, - 64'd50522608463611, - 64'd4844167648166494, - 64'd1362478337710898, 64'd75562184921047, - 64'd48464973598296, - 64'd5505606112695792, - 64'd1283363101544822, 64'd63357707642909, - 64'd46388011318308, - 64'd6127608592846752, - 64'd1204760640672916, 64'd51523776702463, - 64'd44297022280336, - 64'd6710469021378337, - 64'd1126819797494900, 64'd40070597533610, - 64'd42197116997558, - 64'd7254553845721645, - 64'd1049681790049693, 64'd29007126689086, - 64'd40093212685508, - 64'd7760298217955038, - 64'd973480223457806, 64'd18341104403961, - 64'd37990030657636, - 64'd8228202194533767, - 64'd898341117369706, 64'd8079088437795, - 64'd35892094253351, - 64'd8658826953595873, - 64'd824382948694820, - 64'd1773510931011, - 64'd33803727280867, - 64'd9052791037302716, - 64'd751716708883021, - 64'd11212394882350, - 64'd31729052956816, - 64'd9410766626307994, - 64'd680445975029168, - 64'd20234339123830, - 64'd29671993324253, - 64'd9733475853084454, - 64'd610666994071711, - 64'd28837156170178, - 64'd27636269130413, - 64'd10021687160473434, - 64'd542468779358351, - 64'd37019656947158, - 64'd25625400145361, - 64'd10276211711459662, - 64'd475933218855215, - 64'd44781611831252, - 64'd23642705902494, - 64'd10497899855813134, - 64'd411135194280880, - 64'd52123711232892, - 64'd21691306841764, - 64'd10687637658882086, - 64'd348142710452861, - 64'd59047525827604, - 64'd19774125836362, - 64'd10846343497466668, - 64'd287017034141654, - 64'd65555466535783, - 64'd17893890083633, - 64'd10974964727352650, - 64'd227812841736223, - 64'd71650744348217, - 64'd16053133340967}};
	localparam logic signed[63:0] Ffi[0:3][0:79] = '{
		'{- 64'd7789584925020542, 64'd708887221199158, 64'd206702748225345, - 64'd19845819841343, - 64'd7393588604643268, 64'd873085743790186, 64'd189441643064671, - 64'd21110141804839, - 64'd6918639246994867, 64'd1024429359565470, 64'd170276674079435, - 64'd22108944360993, - 64'd6371556198568730, 64'd1161381434685642, 64'd149461551191332, - 64'd22835111110926, - 64'd5759879607888508, 64'd1282597644249564, 64'd127264837936302, - 64'd23284800600437, - 64'd5091771080218742, 64'd1386938313763277, 64'd103966594132111, - 64'd23457435961284, - 64'd4375908801885497, 64'd1473478185138040, 64'd79854941677750, - 64'd23355656937657, - 64'd3621378440744956, 64'd1541513537288885, 64'd55222594523002, - 64'd22985235482842, - 64'd2837561156357778, 64'd1590566623196748, 64'd30363393574268, - 64'd22354956512906, - 64'd2034020064558232, 64'd1620387416998140, 64'd5568886563156, - 64'd21476465781011, - 64'd1220386496487038, 64'd1630952695911008, - 64'd18875008286193, - 64'd20364087183631, - 64'd406247372102465, 64'd1622462512239921, - 64'd42691217575166, - 64'd19034612125145, 64'd398965026813756, 64'd1595334139989243, - 64'd65614571842042, - 64'd17507063846684, 64'd1186079648425665, 64'd1550193608429831, - 64'd87394675671855, - 64'd15802439866300, 64'd1946288454422587, 64'd1487864961015521, - 64'd107798558746626, - 64'd13943435878179, 64'd2671242297735851, 64'd1409357402058381, - 64'd126613080816752, - 64'd11954154617209, 64'd3353139883456778, 64'd1315850515302490, - 64'd143647066875003, - 64'd9859803310541, 64'd3984808899006887, 64'd1208677757771555, - 64'd158733152334642, - 64'd7686383409257, 64'd4559778505553668, 64'd1089308448825112, - 64'd171729321708043, - 64'd5460376320793, 64'd5072342496187033, 64'd959328488094488, - 64'd182520128106280, - 64'd3208428846785},
		'{64'd7789584925020678, - 64'd708887221199165, - 64'd206702748225342, 64'd19845819841342, 64'd7393588604643451, - 64'd873085743790196, - 64'd189441643064668, 64'd21110141804838, 64'd6918639246995094, - 64'd1024429359565484, - 64'd170276674079431, 64'd22108944360992, 64'd6371556198568998, - 64'd1161381434685658, - 64'd149461551191327, 64'd22835111110925, 64'd5759879607888814, - 64'd1282597644249583, - 64'd127264837936296, 64'd23284800600436, 64'd5091771080219080, - 64'd1386938313763298, - 64'd103966594132105, 64'd23457435961283, 64'd4375908801885863, - 64'd1473478185138064, - 64'd79854941677743, 64'd23355656937656, 64'd3621378440745346, - 64'd1541513537288910, - 64'd55222594522994, 64'd22985235482840, 64'd2837561156358186, - 64'd1590566623196775, - 64'd30363393574260, 64'd22354956512905, 64'd2034020064558654, - 64'd1620387416998168, - 64'd5568886563148, 64'd21476465781009, 64'd1220386496487468, - 64'd1630952695911038, 64'd18875008286202, 64'd20364087183629, 64'd406247372102900, - 64'd1622462512239951, 64'd42691217575174, 64'd19034612125143, - 64'd398965026813322, - 64'd1595334139989273, 64'd65614571842050, 64'd17507063846682, - 64'd1186079648425238, - 64'd1550193608429861, 64'd87394675671863, 64'd15802439866299, - 64'd1946288454422172, - 64'd1487864961015550, 64'd107798558746634, 64'd13943435878177, - 64'd2671242297735452, - 64'd1409357402058410, 64'd126613080816760, 64'd11954154617207, - 64'd3353139883456400, - 64'd1315850515302518, 64'd143647066875011, 64'd9859803310540, - 64'd3984808899006532, - 64'd1208677757771581, 64'd158733152334649, 64'd7686383409256, - 64'd4559778505553342, - 64'd1089308448825137, 64'd171729321708049, 64'd5460376320792, - 64'd5072342496186738, - 64'd959328488094511, 64'd182520128106285, 64'd3208428846784},
		'{64'd20410122023596984, - 64'd1087203619517777, 64'd261581401330405, - 64'd19688353631198, 64'd19855845437227768, - 64'd1129165953014674, 64'd260549776479662, - 64'd21497800075813, 64'd19281639300793944, - 64'd1166937977762846, 64'd258996978016206, - 64'd23185429430581, 64'd18689575854732616, - 64'd1200612237457261, 64'd256948048973282, - 64'd24752655664962, 64'd18081679793730520, - 64'd1230286297560720, 64'd254428064696757, - 64'd26201094598827, 64'd17459925861202104, - 64'd1256062325165291, 64'd251462077212791, - 64'd27532552007075, 64'd16826236651983674, - 64'd1278046676369314, 64'd248075061960339, - 64'd28749011807856, 64'd16182480619338714, - 64'd1296349491750649, 64'd244291866905447, - 64'd29852624356494, 64'd15530470282089826, - 64'd1311084300475151, 64'd240137164048391, - 64'd30845694866052, 64'd14871960627433400, - 64'd1322367633538259, 64'd235635403329143, - 64'd31730671974348, 64'd14208647704754270, - 64'd1330318646597064, 64'd230810768931151, - 64'd32510136476076, 64'd13542167405539158, - 64'd1335058752810478, 64'd225687137978284, - 64'd33186790237559, 64'd12874094424288384, - 64'd1336711266066034, 64'd220288041614798, - 64'd33763445310536, 64'd12205941395145922, - 64'd1335401054933668, 64'd214636628453457, - 64'd34243013260277, 64'd11539158198806890, - 64'd1331254207649389, 64'd208755630372409, - 64'd34628494722203, 64'd10875131434119388, - 64'd1324397708395326, 64'd202667330637182, - 64'd34922969200132, 64'd10215184048673250, - 64'd1314959125107046, 64'd196393534320064, - 64'd35129585118164, 64'd9560575122561506, - 64'd1303066309004502, 64'd189955540985356, - 64'd35251550137213, 64'd8912499799410572, - 64'd1288847106009427, 64'd183374119605357, - 64'd35292121746123, 64'd8272089358702066, - 64'd1272429080179444, 64'd176669485668604, - 64'd35254598136332},
		'{- 64'd20410122023597112, 64'd1087203619517783, - 64'd261581401330408, 64'd19688353631199, - 64'd19855845437227944, 64'd1129165953014683, - 64'd260549776479665, 64'd21497800075814, - 64'd19281639300794168, 64'd1166937977762856, - 64'd258996978016210, 64'd23185429430582, - 64'd18689575854732880, 64'd1200612237457274, - 64'd256948048973287, 64'd24752655664963, - 64'd18081679793730820, 64'd1230286297560734, - 64'd254428064696763, 64'd26201094598828, - 64'd17459925861202444, 64'd1256062325165307, - 64'd251462077212797, 64'd27532552007076, - 64'd16826236651984046, 64'd1278046676369332, - 64'd248075061960346, 64'd28749011807857, - 64'd16182480619339120, 64'd1296349491750668, - 64'd244291866905454, 64'd29852624356495, - 64'd15530470282090264, 64'd1311084300475172, - 64'd240137164048399, 64'd30845694866053, - 64'd14871960627433864, 64'd1322367633538281, - 64'd235635403329152, 64'd31730671974350, - 64'd14208647704754760, 64'd1330318646597088, - 64'd230810768931160, 64'd32510136476078, - 64'd13542167405539672, 64'd1335058752810502, - 64'd225687137978293, 64'd33186790237561, - 64'd12874094424288920, 64'd1336711266066060, - 64'd220288041614808, 64'd33763445310538, - 64'd12205941395146478, 64'd1335401054933694, - 64'd214636628453467, 64'd34243013260279, - 64'd11539158198807466, 64'd1331254207649416, - 64'd208755630372419, 64'd34628494722205, - 64'd10875131434119980, 64'd1324397708395354, - 64'd202667330637193, 64'd34922969200134, - 64'd10215184048673856, 64'd1314959125107074, - 64'd196393534320075, 64'd35129585118166, - 64'd9560575122562122, 64'd1303066309004531, - 64'd189955540985367, 64'd35251550137215, - 64'd8912499799411199, 64'd1288847106009456, - 64'd183374119605368, 64'd35292121746125, - 64'd8272089358702702, 64'd1272429080179473, - 64'd176669485668615, 64'd35254598136334}};
	localparam logic signed[63:0] Fbr[0:3][0:79] = '{
		'{- 64'd2678910912348682, 64'd1633669149297615, 64'd134405106412023, - 64'd14489081406757, - 64'd3471761733289509, 64'd1534935316807140, 64'd154547576200402, - 64'd12167341321049, - 64'd4211153497515380, 64'd1420087166233641, 64'd172563932222687, - 64'd9743629047954, - 64'd4889422534499934, 64'd1290723849399400, 64'd188281223922595, - 64'd7247706595933, - 64'd5499740975037776, 64'd1148585763351890, 64'd201556008143343, - 64'd4709673588602, - 64'd6036181793402482, 64'd995532040410431, 64'd212275515540637, - 64'd2159613203878, - 64'd6493772333226378, 64'd833517040657504, 64'd220358442413966, 64'd372755769329, - 64'd6868535890318197, 64'd664566135678268, 64'd225755365061278, 64'd2858416831816, - 64'd7157521071022570, 64'd490751075721102, 64'd228448778179966, 64'd5269379888993, - 64'd7358818790936519, 64'd314165232382821, 64'd228452763163329, 64'd7578988059119, - 64'd7471566924126414, 64'd136899005473061, 64'd225812296327788, 64'd9762203913194, - 64'd7495942755766966, - 64'd38984324020268, 64'd220602211106000, 64'd11795872177577, - 64'd7433143529741519, - 64'd211472022825834, 64'd212925832011491, 64'd13658956252499, - 64'd7285355515665612, - 64'd378624356972050, 64'd202913301681643, 64'd15332746247078, - 64'd7055712145579892, - 64'd538595822537850, 64'd190719625501872, 64'd16801036599608, - 64'd6748241887867779, - 64'd689654930258371, 64'd176522461172683, 64'd18050271736293, - 64'd6367806633571694, - 64'd830202339184127, 64'd160519683075600, 64'd19069658617453, - 64'd5920031467125635, - 64'd958787157130758, 64'd142926753400873, 64'd19851245422781, - 64'd5411226778650929, - 64'd1074121249927379, 64'd123973933701595, 64'd20389966031699, - 64'd4848303747586724, - 64'd1175091427164946, 64'd103903371822373, 64'd20683650356549},
		'{- 64'd2678910912348222, 64'd1633669149297648, 64'd134405106412032, - 64'd14489081406755, - 64'd3471761733289070, 64'd1534935316807172, 64'd154547576200411, - 64'd12167341321048, - 64'd4211153497514966, 64'd1420087166233671, 64'd172563932222695, - 64'd9743629047952, - 64'd4889422534499551, 64'd1290723849399429, 64'd188281223922603, - 64'd7247706595932, - 64'd5499740975037427, 64'd1148585763351916, 64'd201556008143349, - 64'd4709673588600, - 64'd6036181793402171, 64'd995532040410455, 64'd212275515540643, - 64'd2159613203877, - 64'd6493772333226108, 64'd833517040657526, 64'd220358442413972, 64'd372755769330, - 64'd6868535890317968, 64'd664566135678286, 64'd225755365061283, 64'd2858416831817, - 64'd7157521071022387, 64'd490751075721118, 64'd228448778179969, 64'd5269379888994, - 64'd7358818790936382, 64'd314165232382833, 64'd228452763163332, 64'd7578988059119, - 64'd7471566924126326, 64'd136899005473070, 64'd225812296327790, 64'd9762203913194, - 64'd7495942755766923, - 64'd38984324020262, 64'd220602211106001, 64'd11795872177577, - 64'd7433143529741523, - 64'd211472022825831, 64'd212925832011491, 64'd13658956252499, - 64'd7285355515665663, - 64'd378624356972050, 64'd202913301681642, 64'd15332746247078, - 64'd7055712145579987, - 64'd538595822537854, 64'd190719625501870, 64'd16801036599608, - 64'd6748241887867917, - 64'd689654930258378, 64'd176522461172680, 64'd18050271736292, - 64'd6367806633571872, - 64'd830202339184137, 64'd160519683075597, 64'd19069658617452, - 64'd5920031467125852, - 64'd958787157130771, 64'd142926753400869, 64'd19851245422781, - 64'd5411226778651180, - 64'd1074121249927394, 64'd123973933701590, 64'd20389966031698, - 64'd4848303747587006, - 64'd1175091427164964, 64'd103903371822367, 64'd20683650356548},
		'{64'd2621464726625032, - 64'd1601298142322358, - 64'd114277463862052, - 64'd54557765512014, 64'd3402192470904109, - 64'd1521613693668172, - 64'd101035526953527, - 64'd52555428834631, 64'd4143075592769200, - 64'd1441949887694716, - 64'd88125723066021, - 64'd50522608463608, 64'd4844167648167600, - 64'd1362478337710847, - 64'd75562184921028, - 64'd48464973598293, 64'd5505606112696863, - 64'd1283363101544773, - 64'd63357707642890, - 64'd46388011318305, 64'd6127608592847788, - 64'd1204760640672868, - 64'd51523776702445, - 64'd44297022280332, 64'd6710469021379336, - 64'd1126819797494854, - 64'd40070597533593, - 64'd42197116997554, 64'd7254553845722606, - 64'd1049681790049648, - 64'd29007126689070, - 64'd40093212685504, 64'd7760298217955961, - 64'd973480223457764, - 64'd18341104403946, - 64'd37990030657633, 64'd8228202194534652, - 64'd898341117369665, - 64'd8079088437780, - 64'd35892094253348, 64'd8658826953596720, - 64'd824382948694780, 64'd1773510931025, - 64'd33803727280864, 64'd9052791037303526, - 64'd751716708882984, 64'd11212394882364, - 64'd31729052956814, 64'd9410766626308762, - 64'd680445975029133, 64'd20234339123843, - 64'd29671993324251, 64'd9733475853085184, - 64'd610666994071677, 64'd28837156170190, - 64'd27636269130411, 64'd10021687160474126, - 64'd542468779358319, 64'd37019656947170, - 64'd25625400145358, 64'd10276211711460314, - 64'd475933218855185, 64'd44781611831263, - 64'd23642705902492, 64'd10497899855813746, - 64'd411135194280852, 64'd52123711232903, - 64'd21691306841762, 64'd10687637658882664, - 64'd348142710452834, 64'd59047525827614, - 64'd19774125836360, 64'd10846343497467206, - 64'd287017034141629, 64'd65555466535792, - 64'd17893890083631, 64'd10974964727353150, - 64'd227812841736200, 64'd71650744348225, - 64'd16053133340965},
		'{64'd2621464726623828, - 64'd1601298142322414, - 64'd114277463862073, - 64'd54557765512018, 64'd3402192470902937, - 64'd1521613693668227, - 64'd101035526953548, - 64'd52555428834635, 64'd4143075592768060, - 64'd1441949887694769, - 64'd88125723066041, - 64'd50522608463611, 64'd4844167648166494, - 64'd1362478337710898, - 64'd75562184921047, - 64'd48464973598296, 64'd5505606112695792, - 64'd1283363101544822, - 64'd63357707642909, - 64'd46388011318308, 64'd6127608592846752, - 64'd1204760640672916, - 64'd51523776702463, - 64'd44297022280336, 64'd6710469021378337, - 64'd1126819797494900, - 64'd40070597533610, - 64'd42197116997558, 64'd7254553845721645, - 64'd1049681790049693, - 64'd29007126689086, - 64'd40093212685508, 64'd7760298217955038, - 64'd973480223457806, - 64'd18341104403961, - 64'd37990030657636, 64'd8228202194533767, - 64'd898341117369706, - 64'd8079088437795, - 64'd35892094253351, 64'd8658826953595873, - 64'd824382948694820, 64'd1773510931011, - 64'd33803727280867, 64'd9052791037302716, - 64'd751716708883021, 64'd11212394882350, - 64'd31729052956816, 64'd9410766626307994, - 64'd680445975029168, 64'd20234339123830, - 64'd29671993324253, 64'd9733475853084454, - 64'd610666994071711, 64'd28837156170178, - 64'd27636269130413, 64'd10021687160473434, - 64'd542468779358351, 64'd37019656947158, - 64'd25625400145361, 64'd10276211711459662, - 64'd475933218855215, 64'd44781611831252, - 64'd23642705902494, 64'd10497899855813134, - 64'd411135194280880, 64'd52123711232892, - 64'd21691306841764, 64'd10687637658882086, - 64'd348142710452861, 64'd59047525827604, - 64'd19774125836362, 64'd10846343497466668, - 64'd287017034141654, 64'd65555466535783, - 64'd17893890083633, 64'd10974964727352650, - 64'd227812841736223, 64'd71650744348217, - 64'd16053133340967}};
	localparam logic signed[63:0] Fbi[0:3][0:79] = '{
		'{64'd7789584925020542, 64'd708887221199158, - 64'd206702748225345, - 64'd19845819841343, 64'd7393588604643268, 64'd873085743790186, - 64'd189441643064671, - 64'd21110141804839, 64'd6918639246994867, 64'd1024429359565470, - 64'd170276674079435, - 64'd22108944360993, 64'd6371556198568730, 64'd1161381434685642, - 64'd149461551191332, - 64'd22835111110926, 64'd5759879607888508, 64'd1282597644249564, - 64'd127264837936302, - 64'd23284800600437, 64'd5091771080218742, 64'd1386938313763277, - 64'd103966594132111, - 64'd23457435961284, 64'd4375908801885497, 64'd1473478185138040, - 64'd79854941677750, - 64'd23355656937657, 64'd3621378440744956, 64'd1541513537288885, - 64'd55222594523002, - 64'd22985235482842, 64'd2837561156357778, 64'd1590566623196748, - 64'd30363393574268, - 64'd22354956512906, 64'd2034020064558232, 64'd1620387416998140, - 64'd5568886563156, - 64'd21476465781011, 64'd1220386496487038, 64'd1630952695911008, 64'd18875008286193, - 64'd20364087183631, 64'd406247372102465, 64'd1622462512239921, 64'd42691217575166, - 64'd19034612125145, - 64'd398965026813756, 64'd1595334139989243, 64'd65614571842042, - 64'd17507063846684, - 64'd1186079648425665, 64'd1550193608429831, 64'd87394675671855, - 64'd15802439866300, - 64'd1946288454422587, 64'd1487864961015521, 64'd107798558746626, - 64'd13943435878179, - 64'd2671242297735851, 64'd1409357402058381, 64'd126613080816752, - 64'd11954154617209, - 64'd3353139883456778, 64'd1315850515302490, 64'd143647066875003, - 64'd9859803310541, - 64'd3984808899006887, 64'd1208677757771555, 64'd158733152334642, - 64'd7686383409257, - 64'd4559778505553668, 64'd1089308448825112, 64'd171729321708043, - 64'd5460376320793, - 64'd5072342496187033, 64'd959328488094488, 64'd182520128106280, - 64'd3208428846785},
		'{- 64'd7789584925020678, - 64'd708887221199165, 64'd206702748225342, 64'd19845819841342, - 64'd7393588604643451, - 64'd873085743790196, 64'd189441643064668, 64'd21110141804838, - 64'd6918639246995094, - 64'd1024429359565484, 64'd170276674079431, 64'd22108944360992, - 64'd6371556198568998, - 64'd1161381434685658, 64'd149461551191327, 64'd22835111110925, - 64'd5759879607888814, - 64'd1282597644249583, 64'd127264837936296, 64'd23284800600436, - 64'd5091771080219080, - 64'd1386938313763298, 64'd103966594132105, 64'd23457435961283, - 64'd4375908801885863, - 64'd1473478185138064, 64'd79854941677743, 64'd23355656937656, - 64'd3621378440745346, - 64'd1541513537288910, 64'd55222594522994, 64'd22985235482840, - 64'd2837561156358186, - 64'd1590566623196775, 64'd30363393574260, 64'd22354956512905, - 64'd2034020064558654, - 64'd1620387416998168, 64'd5568886563148, 64'd21476465781009, - 64'd1220386496487468, - 64'd1630952695911038, - 64'd18875008286202, 64'd20364087183629, - 64'd406247372102900, - 64'd1622462512239951, - 64'd42691217575174, 64'd19034612125143, 64'd398965026813322, - 64'd1595334139989273, - 64'd65614571842050, 64'd17507063846682, 64'd1186079648425238, - 64'd1550193608429861, - 64'd87394675671863, 64'd15802439866299, 64'd1946288454422172, - 64'd1487864961015550, - 64'd107798558746634, 64'd13943435878177, 64'd2671242297735452, - 64'd1409357402058410, - 64'd126613080816760, 64'd11954154617207, 64'd3353139883456400, - 64'd1315850515302518, - 64'd143647066875011, 64'd9859803310540, 64'd3984808899006532, - 64'd1208677757771581, - 64'd158733152334649, 64'd7686383409256, 64'd4559778505553342, - 64'd1089308448825137, - 64'd171729321708049, 64'd5460376320792, 64'd5072342496186738, - 64'd959328488094511, - 64'd182520128106285, 64'd3208428846784},
		'{- 64'd20410122023596984, - 64'd1087203619517777, - 64'd261581401330405, - 64'd19688353631198, - 64'd19855845437227768, - 64'd1129165953014674, - 64'd260549776479662, - 64'd21497800075813, - 64'd19281639300793944, - 64'd1166937977762846, - 64'd258996978016206, - 64'd23185429430581, - 64'd18689575854732616, - 64'd1200612237457261, - 64'd256948048973282, - 64'd24752655664962, - 64'd18081679793730520, - 64'd1230286297560720, - 64'd254428064696757, - 64'd26201094598827, - 64'd17459925861202104, - 64'd1256062325165291, - 64'd251462077212791, - 64'd27532552007075, - 64'd16826236651983674, - 64'd1278046676369314, - 64'd248075061960339, - 64'd28749011807856, - 64'd16182480619338714, - 64'd1296349491750649, - 64'd244291866905447, - 64'd29852624356494, - 64'd15530470282089826, - 64'd1311084300475151, - 64'd240137164048391, - 64'd30845694866052, - 64'd14871960627433400, - 64'd1322367633538259, - 64'd235635403329143, - 64'd31730671974348, - 64'd14208647704754270, - 64'd1330318646597064, - 64'd230810768931151, - 64'd32510136476076, - 64'd13542167405539158, - 64'd1335058752810478, - 64'd225687137978284, - 64'd33186790237559, - 64'd12874094424288384, - 64'd1336711266066034, - 64'd220288041614798, - 64'd33763445310536, - 64'd12205941395145922, - 64'd1335401054933668, - 64'd214636628453457, - 64'd34243013260277, - 64'd11539158198806890, - 64'd1331254207649389, - 64'd208755630372409, - 64'd34628494722203, - 64'd10875131434119388, - 64'd1324397708395326, - 64'd202667330637182, - 64'd34922969200132, - 64'd10215184048673250, - 64'd1314959125107046, - 64'd196393534320064, - 64'd35129585118164, - 64'd9560575122561506, - 64'd1303066309004502, - 64'd189955540985356, - 64'd35251550137213, - 64'd8912499799410572, - 64'd1288847106009427, - 64'd183374119605357, - 64'd35292121746123, - 64'd8272089358702066, - 64'd1272429080179444, - 64'd176669485668604, - 64'd35254598136332},
		'{64'd20410122023597112, 64'd1087203619517783, 64'd261581401330408, 64'd19688353631199, 64'd19855845437227944, 64'd1129165953014683, 64'd260549776479665, 64'd21497800075814, 64'd19281639300794168, 64'd1166937977762856, 64'd258996978016210, 64'd23185429430582, 64'd18689575854732880, 64'd1200612237457274, 64'd256948048973287, 64'd24752655664963, 64'd18081679793730820, 64'd1230286297560734, 64'd254428064696763, 64'd26201094598828, 64'd17459925861202444, 64'd1256062325165307, 64'd251462077212797, 64'd27532552007076, 64'd16826236651984046, 64'd1278046676369332, 64'd248075061960346, 64'd28749011807857, 64'd16182480619339120, 64'd1296349491750668, 64'd244291866905454, 64'd29852624356495, 64'd15530470282090264, 64'd1311084300475172, 64'd240137164048399, 64'd30845694866053, 64'd14871960627433864, 64'd1322367633538281, 64'd235635403329152, 64'd31730671974350, 64'd14208647704754760, 64'd1330318646597088, 64'd230810768931160, 64'd32510136476078, 64'd13542167405539672, 64'd1335058752810502, 64'd225687137978293, 64'd33186790237561, 64'd12874094424288920, 64'd1336711266066060, 64'd220288041614808, 64'd33763445310538, 64'd12205941395146478, 64'd1335401054933694, 64'd214636628453467, 64'd34243013260279, 64'd11539158198807466, 64'd1331254207649416, 64'd208755630372419, 64'd34628494722205, 64'd10875131434119980, 64'd1324397708395354, 64'd202667330637193, 64'd34922969200134, 64'd10215184048673856, 64'd1314959125107074, 64'd196393534320075, 64'd35129585118166, 64'd9560575122562122, 64'd1303066309004531, 64'd189955540985367, 64'd35251550137215, 64'd8912499799411199, 64'd1288847106009456, 64'd183374119605368, 64'd35292121746125, 64'd8272089358702702, 64'd1272429080179473, 64'd176669485668615, 64'd35254598136334}};
	localparam logic signed[63:0] hf[0:1999] = {64'd7033096503296, - 64'd32897980416, - 64'd10967230464, 64'd63928604, 64'd7000245665792, - 64'd98394423296, - 64'd10337267712, 64'd188110032, 64'd6934845456384, - 64'd162997501952, - 64'd9086782464, 64'd301512896, 64'd6837488844800, - 64'd226124627968, - 64'd7233756672, 64'd397524544, 64'd6709056110592, - 64'd287210536960, - 64'd4804252672, 64'd470098240, 64'd6550703833088, - 64'd345713672192, - 64'd1831931776, 64'd513814560, 64'd6363853881344, - 64'd401122131968, 64'd1642511488, 64'd523933696, 64'd6150172966912, - 64'd452959338496, 64'd5571985920, 64'd496438560, 64'd5911558488064, - 64'd500788854784, 64'd9903706112, 64'd428068320, 64'd5650113888256, - 64'd544219168768, 64'd14579948544, 64'd316342016, 64'd5368126111744, - 64'd582907527168, 64'd19538849792, 64'd159572240, 64'd5068042010624, - 64'd616563212288, 64'd24715249664, - 64'd43130884, 64'd4752438460416, - 64'd644950327296, 64'd30041542656, - 64'd291865696, 64'd4423997194240, - 64'd667889827840, 64'd35448557568, - 64'd585954240, 64'd4085474918400, - 64'd685260537856, 64'd40866439168, - 64'd923966848, 64'd3739673690112, - 64'd697000263680, 64'd46225510400, - 64'd1303755136, 64'd3389412343808, - 64'd703105531904, 64'd51457126400, - 64'd1722493184, 64'd3037497131008, - 64'd703630671872, 64'd56494514176, - 64'd2176726784, 64'd2686692360192, - 64'd698686832640, 64'd61273546752, - 64'd2662427904, 64'd2339693658112, - 64'd688439820288, 64'd65733513216, - 64'd3175056896, 64'd1999099920384, - 64'd673107279872, 64'd69817778176, - 64'd3709628672, 64'd1667389456384, - 64'd652956008448, 64'd73474457600, - 64'd4260784384, 64'd1346895216640, - 64'd628297957376, 64'd76656959488, - 64'd4822863872, 64'd1039784017920, - 64'd599486234624, 64'd79324479488, - 64'd5389984768, 64'd748036685824, - 64'd566910648320, 64'd81442447360, - 64'd5956117504, 64'd473431015424, - 64'd530992660480, 64'd82982838272, - 64'd6515166720, 64'd217527091200, - 64'd492180406272, 64'd83924451328, - 64'd7061048320, - 64'd18344486912, - 64'd450943287296, 64'd84253073408, - 64'd7587765248, - 64'd233092038656, - 64'd407766368256, 64'd83961561088, - 64'd8089484800, - 64'd425869180928, - 64'd363144806400, 64'd83049857024, - 64'd8560607232, - 64'd596078428160, - 64'd317578280960, 64'd81524924416, - 64'd8995835904, - 64'd743372095488, - 64'd271565209600, 64'd79400542208, - 64'd9390236672, - 64'd867650306048, - 64'd225597456384, 64'd76697108480, - 64'd9739302912, - 64'd969056190464, - 64'd180154810368, 64'd73441320960, - 64'd10038998016, - 64'd1047968874496, - 64'd135700045824, 64'd69665783808, - 64'd10285808640, - 64'd1104993583104, - 64'd92673966080, 64'd65408569344, - 64'd10476781568, - 64'd1140949254144, - 64'd51490967552, 64'd60712722432, - 64'd10609551360, - 64'd1156854972416, - 64'd12534914048, 64'd55625695232, - 64'd10682369024, - 64'd1153913061376, 64'd23844581376, 64'd50198769664, - 64'd10694119424, - 64'd1133491388416, 64'd57335398400, 64'd44486422528, - 64'd10644324352, - 64'd1097103966208, 64'd87665672192, 64'd38545653760, - 64'd10533150720, - 64'd1046390308864, 64'd114606071808, 64'd32435316736, - 64'd10361399296, - 64'd983093477376, 64'd137971515392, 64'd26215440384, - 64'd10130492416, - 64'd909037731840, 64'd157622370304, 64'd19946518528, - 64'd9842454528, - 64'd826105724928, 64'd173465124864, 64'd13688829952, - 64'd9499883520, - 64'd736215171072, 64'd185452544000, 64'd7501764608, - 64'd9105917952, - 64'd641296105472, 64'd193583169536, 64'd1443165440, - 64'd8664196096, - 64'd543267749888, 64'd197900484608, - 64'd4431298048, - 64'd8178812416, - 64'd444016885760, 64'd198491455488, - 64'd10068722688, - 64'd7654265856, - 64'd345376227328, 64'd195484614656, - 64'd15419525120, - 64'd7095408640, - 64'd249104269312, 64'd189047783424, - 64'd20437946368, - 64'd6507388928, - 64'd156866412544, 64'd179385237504, - 64'd25082505216, - 64'd5895589888, - 64'd70217392128, 64'd166734675968, - 64'd29316399104, - 64'd5265568768, 64'd9414508544, 64'd151363747840, - 64'd33107843072, - 64'd4622995968, 64'd80741564416, 64'd133566259200, - 64'd36430344192, - 64'd3973589248, 64'd142628683776, 64'd113658347520, - 64'd39262916608, - 64'd3323052544, 64'd194103558144, 64'd91974221824, - 64'd41590218752, - 64'd2677014272, 64'd234364616704, 64'd68861943808, - 64'd43402641408, - 64'd2040966400, 64'd262786842624, 64'd44679032832, - 64'd44696309760, - 64'd1420208256, 64'd278925475840, 64'd19788113920, - 64'd45473042432, - 64'd819790720, 64'd282517438464, - 64'd5447470592, - 64'd45740224512, - 64'd244465792, 64'd273480531968, - 64'd30667960320, - 64'd45510623232, 64'd301360416, 64'd251910750208, - 64'd55521345536, - 64'd44802162688, 64'd813669824, 64'd218077265920, - 64'd79667380224, - 64'd43637624832, 64'd1288869760, 64'd172415664128, - 64'd102781378560, - 64'd42044309504, 64'd1723824640, 64'd115519225856, - 64'd124557795328, - 64'd40053633024, 64'd2115882240, 64'd48128520192, - 64'd144713433088, - 64'd37700722688, 64'd2462894336, - 64'd28880474112, - 64'd162990424064, - 64'd35023921152, 64'd2763230464, - 64'd114509742080, - 64'd179158859776, - 64'd32064319488, 64'd3015787008, - 64'd207653748736, - 64'd193018920960, - 64'd28865234944, 64'd3219988736, - 64'd307115032576, - 64'd204402835456, - 64'd25471664128, 64'd3375784960, - 64'd411620442112, - 64'd213176172544, - 64'd21929756672, 64'd3483641344, - 64'd519838269440, - 64'd219238973440, - 64'd18286260224, 64'd3544522240, - 64'd630395568128, - 64'd222526259200, - 64'd14587981824, 64'd3559872512, - 64'd741895634944, - 64'd223008227328, - 64'd10881244160, 64'd3531590144, - 64'd852935704576, - 64'd220690022400, - 64'd7211374080, 64'd3461996544, - 64'd962124054528, - 64'd215611097088, - 64'd3622200320, 64'd3353801728, - 64'd1068097273856, - 64'd207844130816, - 64'd155578656, 64'd3210066176, - 64'd1169536057344, - 64'd197493669888, 64'd3149049344, 64'd3034159104, - 64'd1265181130752, - 64'd184694308864, 64'd6255063040, 64'd2829713920, - 64'd1353847668736, - 64'd169608675328, 64'd9129030656, 64'd2600581376, - 64'd1434438467584, - 64'd152425005056, 64'd11741032448, 64'd2350781696, - 64'd1505956593664, - 64'd133354577920, 64'd14064936960, 64'd2084455552, - 64'd1567515475968, - 64'd112628752384, 64'd16078633984, 64'd1805813376, - 64'd1618349129728, - 64'd90496016384, 64'd17764208640, 64'd1519086592, - 64'd1657819234304, - 64'd67218747392, 64'd19108071424, 64'd1228478592, - 64'd1685421162496, - 64'd43069902848, 64'd20101029888, 64'd938116672, - 64'd1700789092352, - 64'd18329671680, 64'd20738314240, 64'd652006464, - 64'd1703698104320, 64'd6717959680, 64'd21019545600, 64'd373988160, - 64'd1694065885184, 64'd31788576768, 64'd20948656128, 64'd107695488, - 64'd1671951417344, 64'd56600698880, 64'd20533766144, - 64'd143481952, - 64'd1637553012736, 64'd80879017984, 64'd19787003904, - 64'd376432992, - 64'd1591204642816, 64'd104357543936, 64'd18724286464, - 64'd588355264, - 64'd1533370171392, 64'd126782562304, 64'd17365071872, - 64'd776781440, - 64'd1464636669952, 64'd147915423744, 64'd15732052992, - 64'd939601280, - 64'd1385706160128, 64'd167535099904, 64'd13850836992, - 64'd1075078784, - 64'd1297386569728, 64'd185440518144, 64'd11749591040, - 64'd1181864704, - 64'd1200580722688, 64'd201452535808, 64'd9458661376, - 64'd1259004928, - 64'd1096275197952, 64'd215415816192, 64'd7010174464, - 64'd1305943424, - 64'd985527877632, 64'd227200188416, 64'd4437632000, - 64'd1322520576, - 64'd869455364096, 64'd236701794304, 64'd1775485824, - 64'd1308967168, - 64'd749219348480, 64'd243843940352, - 64'd941283776, - 64'd1265894400, - 64'd626012913664, 64'd248577572864, - 64'd3677590016, - 64'd1194278144, - 64'd501046935552, 64'd250881425408, - 64'd6398656512, - 64'd1095440768, - 64'd375535730688, 64'd250761838592, - 64'd9070423040, - 64'd971028672, - 64'd250683834368, 64'd248252301312, - 64'd11659934720, - 64'd822986240, - 64'd127672295424, 64'd243412647936, - 64'd14135713792, - 64'd653526912, - 64'd7645917696, 64'd236328009728, - 64'd16468104192, - 64'd465101920, 64'd108299083776, 64'd227107389440, - 64'd18629595136, - 64'd260366176, 64'd219126661120, 64'd215882104832, - 64'd20595109888, - 64'd42143052, 64'd323871637504, 64'd202803920896, - 64'd22342254592, 64'd186612704, 64'd421649350656, 64'd188043018240, - 64'd23851552768, 64'd422852640, 64'd511664455680, 64'd171785748480, - 64'd25106614272, 64'd663472896, 64'd593218240512, 64'd154232242176, - 64'd26094284800, 64'd905352320, 64'd665715081216, 64'd135593918464, - 64'd26804754432, 64'd1145390336, 64'd728667193344, 64'd116090904576, - 64'd27231608832, 64'd1380543744, 64'd781698727936, 64'd95949373440, - 64'd27371864064, 64'd1607862400, 64'd824547606528, 64'd75398856704, - 64'd27225939968, 64'd1824522752, 64'd857067028480, 64'd54669598720, - 64'd26797602816, 64'd2027859968, 64'd879224750080, 64'd33989888000, - 64'd26093875200, 64'd2215397376, 64'd891101773824, 64'd13583513600, - 64'd25124898816, 64'd2384873216, 64'd892889333760, - 64'd6332733440, - 64'd23903772672, 64'd2534263552, 64'd884884701184, - 64'd25551407104, - 64'd22446352384, 64'd2661804288, 64'd867486269440, - 64'd43876618240, - 64'd20771020800, 64'd2766007296, 64'd841186934784, - 64'd61126078464, - 64'd18898444288, 64'd2845674240, 64'd806566887424, - 64'd77132947456, - 64'd16851289088, 64'd2899907328, 64'd764285681664, - 64'd91747483648, - 64'd14653930496, 64'd2928114688, 64'd715073060864, - 64'd104838455296, - 64'd12332148736, 64'd2930013696, 64'd659719585792, - 64'd116294311936, - 64'd9912799232, 64'd2905629696, 64'd599066345472, - 64'd126024146944, - 64'd7423496704, 64'd2855291904, 64'd533994668032, - 64'd133958361088, - 64'd4892274176, 64'd2779624704, 64'd465415241728, - 64'd140049088512, - 64'd2347257600, 64'd2679536640, 64'd394257203200, - 64'd144270393344, 64'd183660272, 64'd2556206336, 64'd321457225728, - 64'd146618138624, 64'd2673139712, 64'd2411064576, 64'd247948623872, - 64'd147109675008, 64'd5094700032, 64'd2245774336, 64'd174650785792, - 64'd145783259136, 64'd7423012352, 64'd2062207744, 64'd102458908672, - 64'd142697250816, 64'd9634170880, 64'd1862423296, 64'd32234213376, - 64'd137929080832, 64'd11705949184, 64'd1648637312, - 64'd35205341184, - 64'd131574038528, 64'd13618027520, 64'd1423197824, - 64'd99093577728, - 64'd123743797248, 64'd15352196096, 64'd1188554880, - 64'd158723964928, - 64'd114564939776, 64'd16892532736, 64'd947231424, - 64'd213456617472, - 64'd104177123328, 64'd18225549312, 64'd701792896, - 64'd262724354048, - 64'd92731334656, 64'd19340306432, 64'd454817568, - 64'd306037915648, - 64'd80387866624, 64'd20228497408, 64'd208866800, - 64'd342990127104, - 64'd67314339840, 64'd20884506624, - 64'd33544018, - 64'd373259010048, - 64'd53683642368, 64'd21305427968, - 64'd269973504, - 64'd396609880064, - 64'd39671808000, 64'd21491048448, - 64'd498081024, - 64'd412896460800, - 64'd25455941632, 64'd21443817472, - 64'd715651776, - 64'd422060851200, - 64'd11212149760, 64'd21168769024, - 64'd920620160, - 64'd424132542464, 64'd2886491648, 64'd20673421312, - 64'd1111091072, - 64'd419226353664, 64'd16671883264, 64'd19967651840, - 64'd1285358592, - 64'd407539548160, 64'd29982767104, 64'd19063545856, - 64'd1441922816, - 64'd389347966976, 64'd42666471424, 64'd17975222272, - 64'd1579503232, - 64'd365001244672, 64'd54580543488, 64'd16718628864, - 64'd1697049984, - 64'd334917435392, 64'd65594208256, 64'd15311344640, - 64'd1793752448, - 64'd299576754176, 64'd75589697536, 64'd13772339200, - 64'd1869043840, - 64'd259514777600, 64'd84463378432, 64'd12121732096, - 64'd1922604416, - 64'd215315218432, 64'd92126724096, 64'd10380551168, - 64'd1954360704, - 64'd167602061312, 64'd98507071488, 64'd8570467840, - 64'd1964482176, - 64'd117031575552, 64'd103548190720, 64'd6713540096, - 64'd1953375744, - 64'd64283930624, 64'd107210645504, 64'd4831954432, - 64'd1921676416, - 64'd10054776832, 64'd109471981568, 64'd2947766016, - 64'd1870237312, 64'd44953247744, 64'd110326685696, 64'd1082651264, - 64'd1800114816, 64'd100038934528, 64'd109785948160, - 64'd742337920, - 64'd1712554752, 64'd154510770176, 64'd107877253120, - 64'd2507003392, - 64'd1608973312, 64'd207694921728, 64'd104643788800, - 64'd4192218624, - 64'd1490939392, 64'd258942943232, 64'd100143644672, - 64'd5780130304, - 64'd1360152832, 64'd307638960128, 64'd94448910336, - 64'd7254341120, - 64'd1218423808, 64'd353206403072, 64'd87644585984, - 64'd8600073216, - 64'd1067649472, 64'd395114184704, 64'd79827378176, - 64'd9804311552, - 64'd909791232, 64'd432882253824, 64'd71104356352, - 64'd10855919616, - 64'd746850816, 64'd466086363136, 64'd61591547904, - 64'd11745739776, - 64'd580847104, 64'd494362230784, 64'd51412426752, - 64'd12466658304, - 64'd413792224, 64'd517408784384, 64'd40696356864, - 64'd13013656576, - 64'd247669072, 64'd534990848000, 64'd29576974336, - 64'd13383830528, - 64'd84408840, 64'd546940780544, 64'd18190557184, - 64'd13576387584, 64'd74130096, 64'd553159360512, 64'd6674405888, - 64'd13592614912, 64'd226182256, 64'd553615949824, - 64'd4834780672, - 64'd13435834368, 64'd370093632, 64'd548347740160, - 64'd16202491904, - 64'd13111324672, 64'd504338656, 64'd537458442240, - 64'd27297931264, - 64'd12626223104, 64'd627535488, 64'd521115828224, - 64'd37995479040, - 64'd11989416960, 64'd738459264, 64'd499548880896, - 64'd48176078848, - 64'd11211404288, 64'd836053504, 64'd473044221952, - 64'd57728499712, - 64'd10304146432, 64'd919438912, 64'd441941950464, - 64'd66550517760, - 64'd9280902144, 64'd987920768, 64'd406630694912, - 64'd74549952512, - 64'd8156052992, 64'd1040993088, 64'd367542566912, - 64'd81645584384, - 64'd6944914944, 64'd1078341504, 64'd325147328512, - 64'd87767891968, - 64'd5663543808, 64'd1099843200, 64'd279946461184, - 64'd92859727872, - 64'd4328539136, 64'd1105564672, 64'd232466825216, - 64'd96876699648, - 64'd2956838144, 64'd1095757824, 64'd183254220800, - 64'd99787579392, - 64'd1565513600, 64'd1070853440, 64'd132866760704, - 64'd101574352896, - 64'd171574784, 64'd1031453312, 64'd81868210176, - 64'd102232301568, 64'd1208231424, 64'd978319616, 64'd30821447680, - 64'd101769781248, 64'd2557609472, 64'd912363520, - 64'd19718068224, - 64'd100207943680, 64'd3860898560, 64'd834631680, - 64'd69208547328, - 64'd97580294144, 64'd5103242240, 64'd746291840, - 64'd117127929856, - 64'd93932068864, 64'd6270749696, 64'd648616768, - 64'd162979545088, - 64'd89319563264, 64'd7350639104, 64'd542967744, - 64'd206297481216, - 64'd83809280000, 64'd8331369472, 64'd430777056, - 64'd246651437056, - 64'd77476986880, 64'd9202753536, 64'd313529888, - 64'd283651080192, - 64'd70406725632, 64'd9956050944, 64'd192746128, - 64'd316949954560, - 64'd62689660928, 64'd10584052736, 64'd69961976, - 64'd346248708096, - 64'd54422949888, 64'd11081128960, - 64'd53288364, - 64'd371297878016, - 64'd45708509184, 64'd11443279872, - 64'd175490560, - 64'd391899774976, - 64'd36651757568, 64'd11668144128, - 64'd295167552, - 64'd407910121472, - 64'd27360344064, 64'd11755006976, - 64'd410896192, - 64'd419238739968, - 64'd17942872064, 64'd11704777728, - 64'd521323040, - 64'd425849716736, - 64'd8507630592, 64'd11519951872, - 64'd625179008, - 64'd427760877568, 64'd838650880, 64'd11204558848, - 64'd721292672, - 64'd425042903040, 64'd9992007680, 64'd10764085248, - 64'd808602688, - 64'd417817427968, 64'd18852395008, 64'd10205391872, - 64'd886167872, - 64'd406254944256, 64'd27324768256, 64'd9536608256, - 64'd953176704, - 64'd390571982848, 64'd35320111104, 64'd8767017984, - 64'd1008954368, - 64'd371027836928, 64'd42756349952, 64'd7906931200, - 64'd1052968640, - 64'd347921055744, 64'd49559191552, 64'd6967550976, - 64'd1084833536, - 64'd321585086464, 64'd55662837760, 64'd5960825344, - 64'd1104311424, - 64'd292384145408, 64'd61010624512, 64'd4899297280, - 64'd1111313664, - 64'd260708253696, 64'd65555509248, 64'd3795950592, - 64'd1105899136, - 64'd226968616960, 64'd69260451840, 64'd2664050688, - 64'd1088270976, - 64'd191592300544, 64'd72098676736, 64'd1516986752, - 64'd1058772032, - 64'd155017199616, 64'd74053804032, 64'd368114528, - 64'd1017878592, - 64'd117686788096, 64'd75119886336, - 64'd769398208, - 64'd966192896, - 64'd80044908544, 64'd75301273600, - 64'd1882721152, - 64'd904433792, - 64'd42530721792, 64'd74612400128, - 64'd2959504384, - 64'd833426688, - 64'd5573702144, 64'd73077473280, - 64'd3988013824, - 64'd754092160, 64'd30411114496, 64'd70729965568, - 64'd4957257216, - 64'd667433984, 64'd65027657728, 64'd67612160000, - 64'd5857098752, - 64'd574525888, 64'd97903050752, 64'd63774429184, - 64'd6678363136, - 64'd476498048, 64'd128691486720, 64'd59274575872, - 64'd7412924928, - 64'd374523168, 64'd157077749760, 64'd54177009664, - 64'd8053787136, - 64'd269802144, 64'd182780313600, 64'd48551907328, - 64'd8595142656, - 64'd163549664, 64'd205553975296, 64'd42474287104, - 64'd9032420352, - 64'd56980000, 64'd225192067072, 64'd36023083008, - 64'd9362321408, 64'd48707084, 64'd241528176640, 64'd29280149504, - 64'd9582834688, 64'd152339968, 64'd254437326848, 64'd22329272320, - 64'd9693236224, 64'd252788304, 64'd263836680192, 64'd15255162880, - 64'd9694081024, 64'd348975392, 64'd269685833728, 64'd8142476288, - 64'd9587174400, 64'd439889728, 64'd271986458624, 64'd1074818560, - 64'd9375527936, 64'd524595744, 64'd270781579264, - 64'd5866192896, - 64'd9063308288, 64'd602243328, 64'd266154344448, - 64'd12601840640, - 64'd8655766528, 64'd672076160, 64'd258226323456, - 64'd19057170432, - 64'd8159164928, 64'd733439296, 64'd247155507200, - 64'd25161789440, - 64'd7580680704, 64'd785784512, 64'd233133752320, - 64'd30850611200, - 64'd6928315392, 64'd828675456, 64'd216383995904, - 64'd36064505856, - 64'd6210783744, 64'd861790464, 64'd197157126144, - 64'd40750891008, - 64'd5437403136, 64'd884924608, 64'd175728607232, - 64'd44864233472, - 64'd4617976320, 64'd897990272, 64'd152394776576, - 64'd48366440448, - 64'd3762670080, 64'd901015872, 64'd127469125632, - 64'd51227189248, - 64'd2881891584, 64'd894144000, 64'd101278294016, - 64'd53424144384, - 64'd1986164096, 64'd877627648, 64'd74158080000, - 64'd54943068160, - 64'd1086004096, 64'd851825792, 64'd46449369088, - 64'd55777853440, - 64'd191799792, 64'd817197120, 64'd18494062592, - 64'd55930470400, 64'd686306496, 64'd774293504, - 64'd9368892416, - 64'd55410786304, 64'd1538531200, 64'd723751744, - 64'd36807413760, - 64'd54236319744, 64'd2355556864, 64'd666285184, - 64'd63500029952, - 64'd52431921152, 64'd3128631040, 64'd602673856, - 64'd89139437568, - 64'd50029350912, 64'd3849658368, 64'd533754816, - 64'd113435836416, - 64'd47066787840, 64'd4511283200, 64'd460411168, - 64'd136120008704, - 64'd43588292608, 64'd5106960896, 64'd383561312, - 64'd156946137088, - 64'd39643185152, 64'd5631021568, 64'd304147840, - 64'd175694184448, - 64'd35285385216, 64'd6078718976, 64'd223126112, - 64'd192172146688, - 64'd30572709888, 64'd6446269952, 64'd141453168, - 64'd206217691136, - 64'd25566150656, 64'd6730883584, 64'd60076656, - 64'd217699647488, - 64'd20329084928, 64'd6930774016, - 64'd20075964, - 64'd226518974464, - 64'd14926526464, 64'd7045166592, - 64'd98107728, - 64'd232609366016, - 64'd9424327680, 64'd7074288128, - 64'd173161984, - 64'd235937497088, - 64'd3888407296, 64'd7019345920, - 64'd244431584, - 64'd236502859776, 64'd1616015232, 64'd6882502144, - 64'd311167360, - 64'd234337206272, 64'd7025165824, 64'd6666826240, - 64'd372685728, - 64'd229503696896, 64'd12277432320, 64'd6376248320, - 64'd428375552, - 64'd222095589376, 64'd17314041856, 64'd6015498752, - 64'd477703744, - 64'd212234715136, 64'd22079696896, 64'd5590036992, - 64'd520220320, - 64'd200069513216, 64'd26523152384, 64'd5105980416, - 64'd555562048, - 64'd185772982272, 64'd30597754880, 64'd4570017280, - 64'd583455104, - 64'd169540141056, 64'd34261897216, 64'd3989324800, - 64'd603716864, - 64'd151585505280, 64'd37479415808, 64'd3371473408, - 64'd616256256, - 64'd132140228608, 64'd40219930624, 64'd2724335104, - 64'd621073344, - 64'd111449161728, 64'd42459090944, 64'd2055986048, - 64'd618257728, - 64'd89767772160, 64'd44178755584, 64'd1374610176, - 64'd607985920, - 64'd67359031296, 64'd45367111680, 64'd688401792, - 64'd590518080, - 64'd44490215424, 64'd46018699264, 64'd5471468, - 64'd566193024, - 64'd21429762048, 64'd46134370304, - 64'd666247424, - 64'd535423520, 64'd1555883136, 64'd45721169920, - 64'd1319086976, - 64'd498689888, 64'd24205301760, 64'd44792164352, - 64'd1945729536, - 64'd456533408, 64'd46265061376, 64'd43366166528, - 64'd2539286272, - 64'd409548928, 64'd67492519936, 64'd41467457536, - 64'd3093369600, - 64'd358377120, 64'd87658446848, 64'd39125377024, - 64'd3602159872, - 64'd303696256, 64'd106549485568, 64'd36373929984, - 64'd4060461568, - 64'd246213632, 64'd123970330624, 64'd33251299328, - 64'd4463754240, - 64'd186656976, 64'd139745705984, 64'd29799337984, - 64'd4808232448, - 64'd125765560, 64'd153722093568, 64'd26063024128, - 64'd5090839552, - 64'd64281496, 64'd165769084928, 64'd22089889792, - 64'd5309289472, - 64'd2941044, 64'd175780577280, 64'd17929424896, - 64'd5462078464, 64'd57533836, 64'd183675584512, 64'd13632480256, - 64'd5548493312, 64'd116443600, 64'd189398745088, 64'd9250644992, - 64'd5568603136, 64'd173118880, 64'd192920535040, 64'd4835645952, - 64'd5523246592, 64'd226927712, 64'd194237251584, 64'd438742560, - 64'd5414009344, 64'd277282272, 64'd193370537984, - 64'd3889856000, - 64'd5243192832, 64'd323644960, 64'd190366760960, - 64'd8101555712, - 64'd5013775360, 64'd365533728, 64'd185296093184, - 64'd12149912576, - 64'd4729367040, 64'd402526848, 64'd178251268096, - 64'd15991135232, - 64'd4394157056, 64'd434266688, 64'd169346187264, - 64'd19584544768, - 64'd4012854528, 64'd460462816, 64'd158714167296, - 64'd22892994560, - 64'd3590626816, 64'd480894272, 64'd146506186752, - 64'd25883242496, - 64'd3133030656, 64'd495411008, 64'd132888772608, - 64'd28526272512, - 64'd2645941760, 64'd503934304, 64'd118041862144, - 64'd30797553664, - 64'd2135481216, 64'd506456576, 64'd102156492800, - 64'd32677253120, - 64'd1607940736, 64'd503040352, 64'd85432393728, - 64'd34150387712, - 64'd1069706688, 64'd493816192, 64'd68075581440, - 64'd35206914048, - 64'd527184576, 64'd478980192, 64'd50295820288, - 64'd35841761280, 64'd13275691, 64'd458790528, 64'd32304191488, - 64'd36054810624, 64'd545452224, 64'd433563520, 64'd14310600704, - 64'd35850821632, 64'd1063321216, 64'd403668896, - 64'd3478606336, - 64'd35239272448, 64'd1561123456, 64'd369524608, - 64'd20862973952, - 64'd34234189824, 64'd2033426688, 64'd331591296, - 64'd37650149376, - 64'd32853913600, 64'd2475182848, 64'd290366144, - 64'd53657956352, - 64'd31120795648, 64'd2881780480, 64'd246376544, - 64'd68716351488, - 64'd29060892672, 64'd3249091072, 64'd200173424, - 64'd82669150208, - 64'd26703589376, 64'd3573507840, 64'd152324528, - 64'd95375622144, - 64'd24081211392, 64'd3851980032, 64'd103407576, - 64'd106711851008, - 64'd21228597248, 64'd4082038528, 64'd54003312, - 64'd116571865088, - 64'd18182653952, 64'd4261814272, 64'd4688806, - 64'd124868567040, - 64'd14981902336, 64'd4390051328, - 64'd43969216, - 64'd131534446592, - 64'd11665993728, 64'd4466109440, - 64'd91420760, - 64'd136521965568, - 64'd8275239936, 64'd4489962496, - 64'd137138640, - 64'd139803836416, - 64'd4850135552, 64'd4462188544, - 64'd180624272, - 64'd141372964864, - 64'd1430882688, 64'd4383951872, - 64'd221412864, - 64'd141242171392, 64'd1943064960, 64'd4256981760, - 64'd259078384, - 64'd139443732480, 64'd5233448448, 64'd4083541248, - 64'd293237696, - 64'd136028684288, 64'd8403623936, 64'd3866393344, - 64'd323554464, - 64'd131065856000, 64'd11418961920, 64'd3608760064, - 64'd349742080, - 64'd124640845824, 64'd14247211008, 64'd3314277632, - 64'd371566368, - 64'd116854710272, 64'd16858833920, 64'd2986947328, - 64'd388847200, - 64'd107822514176, 64'd19227299840, 64'd2631084288, - 64'd401459936, - 64'd97671798784, 64'd21329344512, 64'd2251260672, - 64'd409335712, - 64'd86540869632, 64'd23145181184, 64'd1852249216, - 64'd412461504, - 64'd74577018880, 64'd24658677760, 64'd1438965504, - 64'd410879232, - 64'd61934665728, 64'd25857468416, 64'd1016407424, - 64'd404684448, - 64'd48773451776, 64'd26733047808, 64'd589596736, - 64'd394024256, - 64'd35256303616, 64'd27280797696, 64'd163520480, - 64'd379094880, - 64'd21547479040, 64'd27499972608, - 64'd256926192, - 64'd360138432, - 64'd7810651136, 64'd27393648640, - 64'd666995136, - 64'd337439520, 64'd5792974336, 64'd26968619008, - 64'd1062137472, - 64'd311321088, 64'd19106494464, 64'd26235260928, - 64'd1438052992, - 64'd282140192, 64'd31979048960, 64'd25207339008, - 64'd1790736000, - 64'd250283168, 64'd44267466752, 64'd23901808640, - 64'd2116516096, - 64'd216160832, 64'd55837798400, 64'd22338547712, - 64'd2412095488, - 64'd180203184, 64'd66566709248, 64'd20540094464, - 64'd2674580480, - 64'd142854208, 64'd76342730752, 64'd18531325952, - 64'd2901509120, - 64'd104566496, 64'd85067358208, 64'd16339141632, - 64'd3090871296, - 64'd65795828, 64'd92655960064, 64'd13992113152, - 64'd3241124864, - 64'd26995910, 64'd99038543872, 64'd11520123904, - 64'd3351205888, 64'd11386859, 64'd104160296960, 64'd8954007552, - 64'd3420532224, 64'd48918428, 64'd107981996032, 64'd6325167616, - 64'd3449003264, 64'd85181896, 64'd110480179200, 64'd3665207808, - 64'd3436992256, 64'd119782032, 64'd111647170560, 64'd1005561408, - 64'd3385333760, 64'd152349504, 64'd111490867200, - 64'd1622868352, - 64'd3295307008, 64'd182544688, 64'd110034436096, - 64'd4190059008, - 64'd3168613632, 64'd210061120, 64'd107315757056, - 64'd6667201024, - 64'd3007350016, 64'd234628432, 64'd103386734592, - 64'd9027011584, - 64'd2813977088, 64'd256014944, 64'd98312503296, - 64'd11244024832, - 64'd2591285760, 64'd274029632, 64'd92170379264, - 64'd13294855168, - 64'd2342358784, 64'd288523648, 64'd85048827904, - 64'd15158435840, - 64'd2070530560, 64'd299391392, 64'd77046226944, - 64'd16816222208, - 64'd1779343616, 64'd306570976, 64'd68269547520, - 64'd18252363776, - 64'd1472505088, 64'd310044160, 64'd58832982016, - 64'd19453847552, - 64'd1153840384, 64'd309835904, 64'd48856506368, - 64'd20410593280, - 64'd827246976, 64'd306013216, 64'd38464389120, - 64'd21115523072, - 64'd496648352, 64'd298683904, 64'd27783663616, - 64'd21564604416, - 64'd165947968, 64'd287994368, 64'd16942639104, - 64'd21756829696, 64'd161015488, 64'd274127456, 64'd6069367296, - 64'd21694183424, 64'd480511552, 64'd257299680, - 64'd4709823488, - 64'd21381576704, 64'd788959168, 64'd237758064, - 64'd15271768064, - 64'd20826730496, 64'd1082965888, 64'd215776896, - 64'd25497839616, - 64'd20040044544, 64'd1359363712, 64'd191653968, - 64'd35275247616, - 64'd19034429440, 64'd1615242112, 64'd165706880, - 64'd44498239488, - 64'd17825124352, 64'd1847977472, 64'd138268864, - 64'd53069225984, - 64'd16429464576, 64'd2055258368, 64'd109684824, - 64'd60899762176, - 64'd14866663424, 64'd2235107584, 64'd80307000, - 64'd67911417856, - 64'd13157547008, 64'd2385898752, 64'd50490892, - 64'd74036527104, - 64'd11324291072, 64'd2506369792, 64'd20591002, - 64'd79218802688, - 64'd9390139392, 64'd2595631104, - 64'd9043209, - 64'd83413778432, - 64'd7379118592, 64'd2653169920, - 64'd38071296, - 64'd86589120512, - 64'd5315746304, 64'd2678849792, - 64'd66165620, - 64'd88724840448, - 64'd3224739072, 64'd2672905216, - 64'd93014920, - 64'd89813286912, - 64'd1130721792, 64'd2635934208, - 64'd118327656, - 64'd89859039232, 64'd942053824, 64'd2568883456, - 64'd141835040, - 64'd88878645248, 64'd2969985280, 64'd2473032960, - 64'd163293760, - 64'd86900252672, 64'd4930381312, 64'd2349974784, - 64'd182488384, - 64'd83963068416, 64'd6801708544, 64'd2201590016, - 64'd199233408, - 64'd80116711424, 64'd8563822592, 64'd2030020992, - 64'd213374832, - 64'd75420508160, 64'd10198177792, 64'd1837643904, - 64'd224791472, - 64'd69942599680, 64'd11688014848, 64'd1627035520, - 64'd233395808, - 64'd63759036416, 64'd13018524672, 64'd1400941312, - 64'd239134400, - 64'd56952745984, 64'd14176988160, 64'd1162240128, - 64'd241988000, - 64'd49612476416, 64'd15152887808, 64'd913908864, - 64'd241971088, - 64'd41831669760, 64'd15937992704, 64'd658986304, - 64'd239131280, - 64'd33707284480, 64'd16526415872, 64'd400536864, - 64'd233548080, - 64'd25338644480, 64'd16914642944, 64'd141614768, - 64'd225331520, - 64'd16826230784, 64'd17101535232, - 64'd114771248, - 64'd214620368, - 64'd8270504960, 64'd17088299008, - 64'd365691968, - 64'd201579968, 64'd229250672, 64'd16878435328, - 64'd608330368, - 64'd186399968, 64'd8576060928, 64'd16477662208, - 64'd840012160, - 64'd169291648, 64'd16676343808, 64'd15893807104, - 64'd1058234624, - 64'd150485136, 64'd24440932352, 64'd15136688128, - 64'd1260692480, - 64'd130226448, 64'd31786033152, 64'd14217958400, - 64'd1445301760, - 64'd108774312, 64'd38634110976, 64'd13150946304, - 64'd1610219392, - 64'd86397032, 64'd44914671616, 64'd11950475264, - 64'd1753861248, - 64'd63369172, 64'd50564964352, 64'd10632657920, - 64'd1874915968, - 64'd39968276, 64'd55530573824, 64'd9214700544, - 64'd1972355584, - 64'd16471616, 64'd59765919744, 64'd7714673664, - 64'd2045442560, 64'd6847026, 64'd63234625536, 64'd6151298560, - 64'd2093733376, 64'd29720462, 64'd65909788672, 64'd4543711744, - 64'd2117079296, 64'd51891092, 64'd67774132224, 64'd2911243008, - 64'd2115622528, 64'd73113720, 64'd68820041728, 64'd1273183616, - 64'd2089790208, 64'd93158192, 64'd69049499648, - 64'd351433280, - 64'd2040284416, 64'd111811808, 64'd68473896960, - 64'd1944049536, - 64'd1968069376, 64'd128881496, 64'd67113725952, - 64'd3486789120, - 64'd1874356352, 64'd144195728, 64'd64998219776, - 64'd4962652672, - 64'd1760584960, 64'd157606112, 64'd62164844544, - 64'd6355700736, - 64'd1628403200, 64'd168988784, 64'd58658750464, - 64'd7651218944, - 64'd1479644416, 64'd178245392, 64'd54532087808, - 64'd8835868672, - 64'd1316303360, 64'd185303792, 64'd49843318784, - 64'd9897820160, - 64'd1140510208, 64'd190118496, 64'd44656418816, - 64'd10826858496, - 64'd954503680, 64'd192670752, 64'd39040032768, - 64'd11614480384, - 64'd760603392, 64'd192968256, 64'd33066635264, - 64'd12253963264, - 64'd561181504, 64'd191044672, 64'd26811590656, - 64'd12740410368, - 64'd358634592, 64'd186958800, 64'd20352258048, - 64'd13070778368, - 64'd155355344, 64'd180793488, 64'd13767048192, - 64'd13243881472, 64'd46295076, 64'd172654240, 64'd7134508032, - 64'd13260374016, 64'd244013680, 64'd162667648, 64'd532402080, - 64'd13122712576, 64'd435581472, 64'd150979568, - 64'd5963171840, - 64'd12835095552, 64'd618887680, 64'd137753088, - 64'd12278635520, - 64'd12403388416, 64'd791952384, 64'd123166384, - 64'd18343737344, - 64'd11835023360, 64'd952947136, 64'd107410400, - 64'd24092315648, - 64'd11138892800, 64'd1100213760, 64'd90686408, - 64'd29462990848, - 64'd10325217280, 64'd1232280576, 64'd73203528, - 64'd34399793152, - 64'd9405405184, 64'd1347876480, 64'd55176152, - 64'd38852730880, - 64'd8391904768, 64'd1445942016, 64'd36821416, - 64'd42778251264, - 64'd7298036736, 64'd1525638272, 64'd18356602, - 64'd46139658240, - 64'd6137830912, 64'd1586352896, - 64'd3364, - 64'd48907403264, - 64'd4925849088, 64'd1627703296, - 64'd18048354, - 64'd51059314688, - 64'd3677007104, 64'd1649537408, - 64'd35575396, - 64'd52580737024, - 64'd2406398464, 64'd1651931392, - 64'd52390896, - 64'd53464559616, - 64'd1129114624, 64'd1635185152, - 64'd68312728, - 64'd53711183872, 64'd139928944, 64'd1599814784, - 64'd83172152, - 64'd53328396288, 64'd1386162304, 64'd1546543488, - 64'd96815528, - 64'd52331134976, 64'd2595524096, 64'd1476289152, - 64'd109105848, - 64'd50741219328, 64'd3754616064, 64'd1390150784, - 64'd119924056, - 64'd48586973184, 64'd4850846208, 64'd1289392896, - 64'd129170104, - 64'd45902774272, 64'd5872562688, 64'd1175427840, - 64'd136763808, - 64'd42728583168, 64'd6809170432, 64'd1049796992, - 64'd142645424, - 64'd39109353472, 64'd7651239424, 64'd914150976, - 64'd146776032, - 64'd35094458368, 64'd8390590464, 64'd770228544, - 64'd149137584, - 64'd30737025024, 64'd9020372992, 64'd619834944, - 64'd149732832, - 64'd26093264896, 64'd9535118336, 64'd464820192, - 64'd148584864, - 64'd21221765120, 64'd9930782720, 64'd307056544, - 64'd145736576, - 64'd16182777856, 64'd10204768256, 64'd148416656, - 64'd141249808, - 64'd11037487104, 64'd10355931136, - 64'd9248055, - 64'd135204288, - 64'd5847291392, 64'd10384567296, - 64'd164128624, - 64'd127696448, - 64'd673083584, 64'd10292387840, - 64'd314478656, - 64'd118838032, 64'd4425443328, 64'd10082473984, - 64'd458633504, - 64'd108754496, 64'd9390467072, 64'd9759219712, - 64'd595028224, - 64'd97583376, 64'd14166675456, 64'd9328256000, - 64'd722214016, - 64'd85472480, 64'd18701864960, 64'd8796367872, - 64'd838872960, - 64'd72578000, 64'd22947489792, 64'd8171397632, - 64'd943831040, - 64'd59062548, 64'd26859171840, 64'd7462130688, - 64'd1036069504, - 64'd45093212, 64'd30397132800, 64'd6678184448, - 64'd1114734080, - 64'd30839494, 64'd33526589440, 64'd5829879808, - 64'd1179141760, - 64'd16471352, 64'd36218060800, 64'd4928109056, - 64'd1228786048, - 64'd2157196, 64'd38447636480, 64'd3984203008, - 64'd1263340160, 64'd11938022, 64'd40197140480, 64'd3009790464, - 64'd1282657280, 64'd25654662, 64'd41454268416, 64'd2016659712, - 64'd1286769408, 64'd38840152, 64'd42212614144, 64'd1016618176, - 64'd1275884288, 64'd51350640, 64'd42471653376, 64'd21356334, - 64'd1250379776, 64'd63052516, 64'd42236645376, - 64'd957685888, - 64'd1210796416, 64'd73823768, 64'd41518489600, - 64'd1909447296, - 64'd1157828864, 64'd83555224, 64'd40333484032, - 64'd2823367424, - 64'd1092315392, 64'd92151592, 64'd38703067136, - 64'd3689500160, - 64'd1015224960, 64'd99532312, 64'd36653469696, - 64'd4498618368, - 64'd927644736, 64'd105632264, 64'd34215340032, - 64'd5242309120, - 64'd830765056, 64'd110402272, 64'd31423309824, - 64'd5913057792, - 64'd725863872, 64'd113809368, 64'd28315527168, - 64'd6504319488, - 64'd614290688, 64'd115836928, 64'd24933158912, - 64'd7010576896, - 64'd497449664, 64'd116484592, 64'd21319860224, - 64'd7427391488, - 64'd376782464, 64'd115767992, 64'd17521235968, - 64'd7751432704, - 64'd253750912, 64'd113718288, 64'd13584269312, - 64'd7980498432, - 64'd129819680, 64'd110381560, 64'd9556759552, - 64'd8113524224, - 64'd6439408, 64'd105818040, 64'd5486758400, - 64'd8150574080, 64'd114969968, 64'd100101136, 64'd1422006400, - 64'd8092821504, 64'd233035072, 64'd93316416, - 64'd2590614528, - 64'd7942518272, 64'd346444256, 64'd85560352, - 64'd6505608704, - 64'd7702948864, 64'd453961664, 64'd76939064, - 64'd10279368704, - 64'd7378376192, 64'd554440448, 64'd67566928, - 64'd13870651392, - 64'd6973975552, 64'd646834304, 64'd57565096, - 64'd17241012224, - 64'd6495759872, 64'd730208128, 64'd47059976, - 64'd20355205120, - 64'd5950494720, 64'd803746816, 64'd36181704, - 64'd23181537280, - 64'd5345609216, 64'd866762944, 64'd25062552, - 64'd25692176384, - 64'd4689098240, 64'd918702144, 64'd13835381, - 64'd27863408640, - 64'd3989420544, 64'd959147840, 64'd2632072, - 64'd29675841536, - 64'd3255392000, 64'd987823232, - 64'd8417969, - 64'd31114557440, - 64'd2496078848, 64'd1004592512, - 64'd19189274, - 64'd32169211904, - 64'd1720688896, 64'd1009460096, - 64'd29561700, - 64'd32834078720, - 64'd938460864, 64'd1002568000, - 64'd39421732, - 64'd33108035584, - 64'd158558640, 64'd984192000, - 64'd48663680, - 64'd32994498560, 64'd610034432, 64'd954736192, - 64'd57190776};
	localparam logic signed[63:0] hb[0:1999] = {64'd7033096503296, 64'd32897980416, - 64'd10967230464, - 64'd63928604, 64'd7000245665792, 64'd98394423296, - 64'd10337267712, - 64'd188110032, 64'd6934845456384, 64'd162997501952, - 64'd9086782464, - 64'd301512896, 64'd6837488844800, 64'd226124627968, - 64'd7233756672, - 64'd397524544, 64'd6709056110592, 64'd287210536960, - 64'd4804252672, - 64'd470098240, 64'd6550703833088, 64'd345713672192, - 64'd1831931776, - 64'd513814560, 64'd6363853881344, 64'd401122131968, 64'd1642511488, - 64'd523933696, 64'd6150172966912, 64'd452959338496, 64'd5571985920, - 64'd496438560, 64'd5911558488064, 64'd500788854784, 64'd9903706112, - 64'd428068320, 64'd5650113888256, 64'd544219168768, 64'd14579948544, - 64'd316342016, 64'd5368126111744, 64'd582907527168, 64'd19538849792, - 64'd159572240, 64'd5068042010624, 64'd616563212288, 64'd24715249664, 64'd43130884, 64'd4752438460416, 64'd644950327296, 64'd30041542656, 64'd291865696, 64'd4423997194240, 64'd667889827840, 64'd35448557568, 64'd585954240, 64'd4085474918400, 64'd685260537856, 64'd40866439168, 64'd923966848, 64'd3739673690112, 64'd697000263680, 64'd46225510400, 64'd1303755136, 64'd3389412343808, 64'd703105531904, 64'd51457126400, 64'd1722493184, 64'd3037497131008, 64'd703630671872, 64'd56494514176, 64'd2176726784, 64'd2686692360192, 64'd698686832640, 64'd61273546752, 64'd2662427904, 64'd2339693658112, 64'd688439820288, 64'd65733513216, 64'd3175056896, 64'd1999099920384, 64'd673107279872, 64'd69817778176, 64'd3709628672, 64'd1667389456384, 64'd652956008448, 64'd73474457600, 64'd4260784384, 64'd1346895216640, 64'd628297957376, 64'd76656959488, 64'd4822863872, 64'd1039784017920, 64'd599486234624, 64'd79324479488, 64'd5389984768, 64'd748036685824, 64'd566910648320, 64'd81442447360, 64'd5956117504, 64'd473431015424, 64'd530992660480, 64'd82982838272, 64'd6515166720, 64'd217527091200, 64'd492180406272, 64'd83924451328, 64'd7061048320, - 64'd18344486912, 64'd450943287296, 64'd84253073408, 64'd7587765248, - 64'd233092038656, 64'd407766368256, 64'd83961561088, 64'd8089484800, - 64'd425869180928, 64'd363144806400, 64'd83049857024, 64'd8560607232, - 64'd596078428160, 64'd317578280960, 64'd81524924416, 64'd8995835904, - 64'd743372095488, 64'd271565209600, 64'd79400542208, 64'd9390236672, - 64'd867650306048, 64'd225597456384, 64'd76697108480, 64'd9739302912, - 64'd969056190464, 64'd180154810368, 64'd73441320960, 64'd10038998016, - 64'd1047968874496, 64'd135700045824, 64'd69665783808, 64'd10285808640, - 64'd1104993583104, 64'd92673966080, 64'd65408569344, 64'd10476781568, - 64'd1140949254144, 64'd51490967552, 64'd60712722432, 64'd10609551360, - 64'd1156854972416, 64'd12534914048, 64'd55625695232, 64'd10682369024, - 64'd1153913061376, - 64'd23844581376, 64'd50198769664, 64'd10694119424, - 64'd1133491388416, - 64'd57335398400, 64'd44486422528, 64'd10644324352, - 64'd1097103966208, - 64'd87665672192, 64'd38545653760, 64'd10533150720, - 64'd1046390308864, - 64'd114606071808, 64'd32435316736, 64'd10361399296, - 64'd983093477376, - 64'd137971515392, 64'd26215440384, 64'd10130492416, - 64'd909037731840, - 64'd157622370304, 64'd19946518528, 64'd9842454528, - 64'd826105724928, - 64'd173465124864, 64'd13688829952, 64'd9499883520, - 64'd736215171072, - 64'd185452544000, 64'd7501764608, 64'd9105917952, - 64'd641296105472, - 64'd193583169536, 64'd1443165440, 64'd8664196096, - 64'd543267749888, - 64'd197900484608, - 64'd4431298048, 64'd8178812416, - 64'd444016885760, - 64'd198491455488, - 64'd10068722688, 64'd7654265856, - 64'd345376227328, - 64'd195484614656, - 64'd15419525120, 64'd7095408640, - 64'd249104269312, - 64'd189047783424, - 64'd20437946368, 64'd6507388928, - 64'd156866412544, - 64'd179385237504, - 64'd25082505216, 64'd5895589888, - 64'd70217392128, - 64'd166734675968, - 64'd29316399104, 64'd5265568768, 64'd9414508544, - 64'd151363747840, - 64'd33107843072, 64'd4622995968, 64'd80741564416, - 64'd133566259200, - 64'd36430344192, 64'd3973589248, 64'd142628683776, - 64'd113658347520, - 64'd39262916608, 64'd3323052544, 64'd194103558144, - 64'd91974221824, - 64'd41590218752, 64'd2677014272, 64'd234364616704, - 64'd68861943808, - 64'd43402641408, 64'd2040966400, 64'd262786842624, - 64'd44679032832, - 64'd44696309760, 64'd1420208256, 64'd278925475840, - 64'd19788113920, - 64'd45473042432, 64'd819790720, 64'd282517438464, 64'd5447470592, - 64'd45740224512, 64'd244465792, 64'd273480531968, 64'd30667960320, - 64'd45510623232, - 64'd301360416, 64'd251910750208, 64'd55521345536, - 64'd44802162688, - 64'd813669824, 64'd218077265920, 64'd79667380224, - 64'd43637624832, - 64'd1288869760, 64'd172415664128, 64'd102781378560, - 64'd42044309504, - 64'd1723824640, 64'd115519225856, 64'd124557795328, - 64'd40053633024, - 64'd2115882240, 64'd48128520192, 64'd144713433088, - 64'd37700722688, - 64'd2462894336, - 64'd28880474112, 64'd162990424064, - 64'd35023921152, - 64'd2763230464, - 64'd114509742080, 64'd179158859776, - 64'd32064319488, - 64'd3015787008, - 64'd207653748736, 64'd193018920960, - 64'd28865234944, - 64'd3219988736, - 64'd307115032576, 64'd204402835456, - 64'd25471664128, - 64'd3375784960, - 64'd411620442112, 64'd213176172544, - 64'd21929756672, - 64'd3483641344, - 64'd519838269440, 64'd219238973440, - 64'd18286260224, - 64'd3544522240, - 64'd630395568128, 64'd222526259200, - 64'd14587981824, - 64'd3559872512, - 64'd741895634944, 64'd223008227328, - 64'd10881244160, - 64'd3531590144, - 64'd852935704576, 64'd220690022400, - 64'd7211374080, - 64'd3461996544, - 64'd962124054528, 64'd215611097088, - 64'd3622200320, - 64'd3353801728, - 64'd1068097273856, 64'd207844130816, - 64'd155578656, - 64'd3210066176, - 64'd1169536057344, 64'd197493669888, 64'd3149049344, - 64'd3034159104, - 64'd1265181130752, 64'd184694308864, 64'd6255063040, - 64'd2829713920, - 64'd1353847668736, 64'd169608675328, 64'd9129030656, - 64'd2600581376, - 64'd1434438467584, 64'd152425005056, 64'd11741032448, - 64'd2350781696, - 64'd1505956593664, 64'd133354577920, 64'd14064936960, - 64'd2084455552, - 64'd1567515475968, 64'd112628752384, 64'd16078633984, - 64'd1805813376, - 64'd1618349129728, 64'd90496016384, 64'd17764208640, - 64'd1519086592, - 64'd1657819234304, 64'd67218747392, 64'd19108071424, - 64'd1228478592, - 64'd1685421162496, 64'd43069902848, 64'd20101029888, - 64'd938116672, - 64'd1700789092352, 64'd18329671680, 64'd20738314240, - 64'd652006464, - 64'd1703698104320, - 64'd6717959680, 64'd21019545600, - 64'd373988160, - 64'd1694065885184, - 64'd31788576768, 64'd20948656128, - 64'd107695488, - 64'd1671951417344, - 64'd56600698880, 64'd20533766144, 64'd143481952, - 64'd1637553012736, - 64'd80879017984, 64'd19787003904, 64'd376432992, - 64'd1591204642816, - 64'd104357543936, 64'd18724286464, 64'd588355264, - 64'd1533370171392, - 64'd126782562304, 64'd17365071872, 64'd776781440, - 64'd1464636669952, - 64'd147915423744, 64'd15732052992, 64'd939601280, - 64'd1385706160128, - 64'd167535099904, 64'd13850836992, 64'd1075078784, - 64'd1297386569728, - 64'd185440518144, 64'd11749591040, 64'd1181864704, - 64'd1200580722688, - 64'd201452535808, 64'd9458661376, 64'd1259004928, - 64'd1096275197952, - 64'd215415816192, 64'd7010174464, 64'd1305943424, - 64'd985527877632, - 64'd227200188416, 64'd4437632000, 64'd1322520576, - 64'd869455364096, - 64'd236701794304, 64'd1775485824, 64'd1308967168, - 64'd749219348480, - 64'd243843940352, - 64'd941283776, 64'd1265894400, - 64'd626012913664, - 64'd248577572864, - 64'd3677590016, 64'd1194278144, - 64'd501046935552, - 64'd250881425408, - 64'd6398656512, 64'd1095440768, - 64'd375535730688, - 64'd250761838592, - 64'd9070423040, 64'd971028672, - 64'd250683834368, - 64'd248252301312, - 64'd11659934720, 64'd822986240, - 64'd127672295424, - 64'd243412647936, - 64'd14135713792, 64'd653526912, - 64'd7645917696, - 64'd236328009728, - 64'd16468104192, 64'd465101920, 64'd108299083776, - 64'd227107389440, - 64'd18629595136, 64'd260366176, 64'd219126661120, - 64'd215882104832, - 64'd20595109888, 64'd42143052, 64'd323871637504, - 64'd202803920896, - 64'd22342254592, - 64'd186612704, 64'd421649350656, - 64'd188043018240, - 64'd23851552768, - 64'd422852640, 64'd511664455680, - 64'd171785748480, - 64'd25106614272, - 64'd663472896, 64'd593218240512, - 64'd154232242176, - 64'd26094284800, - 64'd905352320, 64'd665715081216, - 64'd135593918464, - 64'd26804754432, - 64'd1145390336, 64'd728667193344, - 64'd116090904576, - 64'd27231608832, - 64'd1380543744, 64'd781698727936, - 64'd95949373440, - 64'd27371864064, - 64'd1607862400, 64'd824547606528, - 64'd75398856704, - 64'd27225939968, - 64'd1824522752, 64'd857067028480, - 64'd54669598720, - 64'd26797602816, - 64'd2027859968, 64'd879224750080, - 64'd33989888000, - 64'd26093875200, - 64'd2215397376, 64'd891101773824, - 64'd13583513600, - 64'd25124898816, - 64'd2384873216, 64'd892889333760, 64'd6332733440, - 64'd23903772672, - 64'd2534263552, 64'd884884701184, 64'd25551407104, - 64'd22446352384, - 64'd2661804288, 64'd867486269440, 64'd43876618240, - 64'd20771020800, - 64'd2766007296, 64'd841186934784, 64'd61126078464, - 64'd18898444288, - 64'd2845674240, 64'd806566887424, 64'd77132947456, - 64'd16851289088, - 64'd2899907328, 64'd764285681664, 64'd91747483648, - 64'd14653930496, - 64'd2928114688, 64'd715073060864, 64'd104838455296, - 64'd12332148736, - 64'd2930013696, 64'd659719585792, 64'd116294311936, - 64'd9912799232, - 64'd2905629696, 64'd599066345472, 64'd126024146944, - 64'd7423496704, - 64'd2855291904, 64'd533994668032, 64'd133958361088, - 64'd4892274176, - 64'd2779624704, 64'd465415241728, 64'd140049088512, - 64'd2347257600, - 64'd2679536640, 64'd394257203200, 64'd144270393344, 64'd183660272, - 64'd2556206336, 64'd321457225728, 64'd146618138624, 64'd2673139712, - 64'd2411064576, 64'd247948623872, 64'd147109675008, 64'd5094700032, - 64'd2245774336, 64'd174650785792, 64'd145783259136, 64'd7423012352, - 64'd2062207744, 64'd102458908672, 64'd142697250816, 64'd9634170880, - 64'd1862423296, 64'd32234213376, 64'd137929080832, 64'd11705949184, - 64'd1648637312, - 64'd35205341184, 64'd131574038528, 64'd13618027520, - 64'd1423197824, - 64'd99093577728, 64'd123743797248, 64'd15352196096, - 64'd1188554880, - 64'd158723964928, 64'd114564939776, 64'd16892532736, - 64'd947231424, - 64'd213456617472, 64'd104177123328, 64'd18225549312, - 64'd701792896, - 64'd262724354048, 64'd92731334656, 64'd19340306432, - 64'd454817568, - 64'd306037915648, 64'd80387866624, 64'd20228497408, - 64'd208866800, - 64'd342990127104, 64'd67314339840, 64'd20884506624, 64'd33544018, - 64'd373259010048, 64'd53683642368, 64'd21305427968, 64'd269973504, - 64'd396609880064, 64'd39671808000, 64'd21491048448, 64'd498081024, - 64'd412896460800, 64'd25455941632, 64'd21443817472, 64'd715651776, - 64'd422060851200, 64'd11212149760, 64'd21168769024, 64'd920620160, - 64'd424132542464, - 64'd2886491648, 64'd20673421312, 64'd1111091072, - 64'd419226353664, - 64'd16671883264, 64'd19967651840, 64'd1285358592, - 64'd407539548160, - 64'd29982767104, 64'd19063545856, 64'd1441922816, - 64'd389347966976, - 64'd42666471424, 64'd17975222272, 64'd1579503232, - 64'd365001244672, - 64'd54580543488, 64'd16718628864, 64'd1697049984, - 64'd334917435392, - 64'd65594208256, 64'd15311344640, 64'd1793752448, - 64'd299576754176, - 64'd75589697536, 64'd13772339200, 64'd1869043840, - 64'd259514777600, - 64'd84463378432, 64'd12121732096, 64'd1922604416, - 64'd215315218432, - 64'd92126724096, 64'd10380551168, 64'd1954360704, - 64'd167602061312, - 64'd98507071488, 64'd8570467840, 64'd1964482176, - 64'd117031575552, - 64'd103548190720, 64'd6713540096, 64'd1953375744, - 64'd64283930624, - 64'd107210645504, 64'd4831954432, 64'd1921676416, - 64'd10054776832, - 64'd109471981568, 64'd2947766016, 64'd1870237312, 64'd44953247744, - 64'd110326685696, 64'd1082651264, 64'd1800114816, 64'd100038934528, - 64'd109785948160, - 64'd742337920, 64'd1712554752, 64'd154510770176, - 64'd107877253120, - 64'd2507003392, 64'd1608973312, 64'd207694921728, - 64'd104643788800, - 64'd4192218624, 64'd1490939392, 64'd258942943232, - 64'd100143644672, - 64'd5780130304, 64'd1360152832, 64'd307638960128, - 64'd94448910336, - 64'd7254341120, 64'd1218423808, 64'd353206403072, - 64'd87644585984, - 64'd8600073216, 64'd1067649472, 64'd395114184704, - 64'd79827378176, - 64'd9804311552, 64'd909791232, 64'd432882253824, - 64'd71104356352, - 64'd10855919616, 64'd746850816, 64'd466086363136, - 64'd61591547904, - 64'd11745739776, 64'd580847104, 64'd494362230784, - 64'd51412426752, - 64'd12466658304, 64'd413792224, 64'd517408784384, - 64'd40696356864, - 64'd13013656576, 64'd247669072, 64'd534990848000, - 64'd29576974336, - 64'd13383830528, 64'd84408840, 64'd546940780544, - 64'd18190557184, - 64'd13576387584, - 64'd74130096, 64'd553159360512, - 64'd6674405888, - 64'd13592614912, - 64'd226182256, 64'd553615949824, 64'd4834780672, - 64'd13435834368, - 64'd370093632, 64'd548347740160, 64'd16202491904, - 64'd13111324672, - 64'd504338656, 64'd537458442240, 64'd27297931264, - 64'd12626223104, - 64'd627535488, 64'd521115828224, 64'd37995479040, - 64'd11989416960, - 64'd738459264, 64'd499548880896, 64'd48176078848, - 64'd11211404288, - 64'd836053504, 64'd473044221952, 64'd57728499712, - 64'd10304146432, - 64'd919438912, 64'd441941950464, 64'd66550517760, - 64'd9280902144, - 64'd987920768, 64'd406630694912, 64'd74549952512, - 64'd8156052992, - 64'd1040993088, 64'd367542566912, 64'd81645584384, - 64'd6944914944, - 64'd1078341504, 64'd325147328512, 64'd87767891968, - 64'd5663543808, - 64'd1099843200, 64'd279946461184, 64'd92859727872, - 64'd4328539136, - 64'd1105564672, 64'd232466825216, 64'd96876699648, - 64'd2956838144, - 64'd1095757824, 64'd183254220800, 64'd99787579392, - 64'd1565513600, - 64'd1070853440, 64'd132866760704, 64'd101574352896, - 64'd171574784, - 64'd1031453312, 64'd81868210176, 64'd102232301568, 64'd1208231424, - 64'd978319616, 64'd30821447680, 64'd101769781248, 64'd2557609472, - 64'd912363520, - 64'd19718068224, 64'd100207943680, 64'd3860898560, - 64'd834631680, - 64'd69208547328, 64'd97580294144, 64'd5103242240, - 64'd746291840, - 64'd117127929856, 64'd93932068864, 64'd6270749696, - 64'd648616768, - 64'd162979545088, 64'd89319563264, 64'd7350639104, - 64'd542967744, - 64'd206297481216, 64'd83809280000, 64'd8331369472, - 64'd430777056, - 64'd246651437056, 64'd77476986880, 64'd9202753536, - 64'd313529888, - 64'd283651080192, 64'd70406725632, 64'd9956050944, - 64'd192746128, - 64'd316949954560, 64'd62689660928, 64'd10584052736, - 64'd69961976, - 64'd346248708096, 64'd54422949888, 64'd11081128960, 64'd53288364, - 64'd371297878016, 64'd45708509184, 64'd11443279872, 64'd175490560, - 64'd391899774976, 64'd36651757568, 64'd11668144128, 64'd295167552, - 64'd407910121472, 64'd27360344064, 64'd11755006976, 64'd410896192, - 64'd419238739968, 64'd17942872064, 64'd11704777728, 64'd521323040, - 64'd425849716736, 64'd8507630592, 64'd11519951872, 64'd625179008, - 64'd427760877568, - 64'd838650880, 64'd11204558848, 64'd721292672, - 64'd425042903040, - 64'd9992007680, 64'd10764085248, 64'd808602688, - 64'd417817427968, - 64'd18852395008, 64'd10205391872, 64'd886167872, - 64'd406254944256, - 64'd27324768256, 64'd9536608256, 64'd953176704, - 64'd390571982848, - 64'd35320111104, 64'd8767017984, 64'd1008954368, - 64'd371027836928, - 64'd42756349952, 64'd7906931200, 64'd1052968640, - 64'd347921055744, - 64'd49559191552, 64'd6967550976, 64'd1084833536, - 64'd321585086464, - 64'd55662837760, 64'd5960825344, 64'd1104311424, - 64'd292384145408, - 64'd61010624512, 64'd4899297280, 64'd1111313664, - 64'd260708253696, - 64'd65555509248, 64'd3795950592, 64'd1105899136, - 64'd226968616960, - 64'd69260451840, 64'd2664050688, 64'd1088270976, - 64'd191592300544, - 64'd72098676736, 64'd1516986752, 64'd1058772032, - 64'd155017199616, - 64'd74053804032, 64'd368114528, 64'd1017878592, - 64'd117686788096, - 64'd75119886336, - 64'd769398208, 64'd966192896, - 64'd80044908544, - 64'd75301273600, - 64'd1882721152, 64'd904433792, - 64'd42530721792, - 64'd74612400128, - 64'd2959504384, 64'd833426688, - 64'd5573702144, - 64'd73077473280, - 64'd3988013824, 64'd754092160, 64'd30411114496, - 64'd70729965568, - 64'd4957257216, 64'd667433984, 64'd65027657728, - 64'd67612160000, - 64'd5857098752, 64'd574525888, 64'd97903050752, - 64'd63774429184, - 64'd6678363136, 64'd476498048, 64'd128691486720, - 64'd59274575872, - 64'd7412924928, 64'd374523168, 64'd157077749760, - 64'd54177009664, - 64'd8053787136, 64'd269802144, 64'd182780313600, - 64'd48551907328, - 64'd8595142656, 64'd163549664, 64'd205553975296, - 64'd42474287104, - 64'd9032420352, 64'd56980000, 64'd225192067072, - 64'd36023083008, - 64'd9362321408, - 64'd48707084, 64'd241528176640, - 64'd29280149504, - 64'd9582834688, - 64'd152339968, 64'd254437326848, - 64'd22329272320, - 64'd9693236224, - 64'd252788304, 64'd263836680192, - 64'd15255162880, - 64'd9694081024, - 64'd348975392, 64'd269685833728, - 64'd8142476288, - 64'd9587174400, - 64'd439889728, 64'd271986458624, - 64'd1074818560, - 64'd9375527936, - 64'd524595744, 64'd270781579264, 64'd5866192896, - 64'd9063308288, - 64'd602243328, 64'd266154344448, 64'd12601840640, - 64'd8655766528, - 64'd672076160, 64'd258226323456, 64'd19057170432, - 64'd8159164928, - 64'd733439296, 64'd247155507200, 64'd25161789440, - 64'd7580680704, - 64'd785784512, 64'd233133752320, 64'd30850611200, - 64'd6928315392, - 64'd828675456, 64'd216383995904, 64'd36064505856, - 64'd6210783744, - 64'd861790464, 64'd197157126144, 64'd40750891008, - 64'd5437403136, - 64'd884924608, 64'd175728607232, 64'd44864233472, - 64'd4617976320, - 64'd897990272, 64'd152394776576, 64'd48366440448, - 64'd3762670080, - 64'd901015872, 64'd127469125632, 64'd51227189248, - 64'd2881891584, - 64'd894144000, 64'd101278294016, 64'd53424144384, - 64'd1986164096, - 64'd877627648, 64'd74158080000, 64'd54943068160, - 64'd1086004096, - 64'd851825792, 64'd46449369088, 64'd55777853440, - 64'd191799792, - 64'd817197120, 64'd18494062592, 64'd55930470400, 64'd686306496, - 64'd774293504, - 64'd9368892416, 64'd55410786304, 64'd1538531200, - 64'd723751744, - 64'd36807413760, 64'd54236319744, 64'd2355556864, - 64'd666285184, - 64'd63500029952, 64'd52431921152, 64'd3128631040, - 64'd602673856, - 64'd89139437568, 64'd50029350912, 64'd3849658368, - 64'd533754816, - 64'd113435836416, 64'd47066787840, 64'd4511283200, - 64'd460411168, - 64'd136120008704, 64'd43588292608, 64'd5106960896, - 64'd383561312, - 64'd156946137088, 64'd39643185152, 64'd5631021568, - 64'd304147840, - 64'd175694184448, 64'd35285385216, 64'd6078718976, - 64'd223126112, - 64'd192172146688, 64'd30572709888, 64'd6446269952, - 64'd141453168, - 64'd206217691136, 64'd25566150656, 64'd6730883584, - 64'd60076656, - 64'd217699647488, 64'd20329084928, 64'd6930774016, 64'd20075964, - 64'd226518974464, 64'd14926526464, 64'd7045166592, 64'd98107728, - 64'd232609366016, 64'd9424327680, 64'd7074288128, 64'd173161984, - 64'd235937497088, 64'd3888407296, 64'd7019345920, 64'd244431584, - 64'd236502859776, - 64'd1616015232, 64'd6882502144, 64'd311167360, - 64'd234337206272, - 64'd7025165824, 64'd6666826240, 64'd372685728, - 64'd229503696896, - 64'd12277432320, 64'd6376248320, 64'd428375552, - 64'd222095589376, - 64'd17314041856, 64'd6015498752, 64'd477703744, - 64'd212234715136, - 64'd22079696896, 64'd5590036992, 64'd520220320, - 64'd200069513216, - 64'd26523152384, 64'd5105980416, 64'd555562048, - 64'd185772982272, - 64'd30597754880, 64'd4570017280, 64'd583455104, - 64'd169540141056, - 64'd34261897216, 64'd3989324800, 64'd603716864, - 64'd151585505280, - 64'd37479415808, 64'd3371473408, 64'd616256256, - 64'd132140228608, - 64'd40219930624, 64'd2724335104, 64'd621073344, - 64'd111449161728, - 64'd42459090944, 64'd2055986048, 64'd618257728, - 64'd89767772160, - 64'd44178755584, 64'd1374610176, 64'd607985920, - 64'd67359031296, - 64'd45367111680, 64'd688401792, 64'd590518080, - 64'd44490215424, - 64'd46018699264, 64'd5471468, 64'd566193024, - 64'd21429762048, - 64'd46134370304, - 64'd666247424, 64'd535423520, 64'd1555883136, - 64'd45721169920, - 64'd1319086976, 64'd498689888, 64'd24205301760, - 64'd44792164352, - 64'd1945729536, 64'd456533408, 64'd46265061376, - 64'd43366166528, - 64'd2539286272, 64'd409548928, 64'd67492519936, - 64'd41467457536, - 64'd3093369600, 64'd358377120, 64'd87658446848, - 64'd39125377024, - 64'd3602159872, 64'd303696256, 64'd106549485568, - 64'd36373929984, - 64'd4060461568, 64'd246213632, 64'd123970330624, - 64'd33251299328, - 64'd4463754240, 64'd186656976, 64'd139745705984, - 64'd29799337984, - 64'd4808232448, 64'd125765560, 64'd153722093568, - 64'd26063024128, - 64'd5090839552, 64'd64281496, 64'd165769084928, - 64'd22089889792, - 64'd5309289472, 64'd2941044, 64'd175780577280, - 64'd17929424896, - 64'd5462078464, - 64'd57533836, 64'd183675584512, - 64'd13632480256, - 64'd5548493312, - 64'd116443600, 64'd189398745088, - 64'd9250644992, - 64'd5568603136, - 64'd173118880, 64'd192920535040, - 64'd4835645952, - 64'd5523246592, - 64'd226927712, 64'd194237251584, - 64'd438742560, - 64'd5414009344, - 64'd277282272, 64'd193370537984, 64'd3889856000, - 64'd5243192832, - 64'd323644960, 64'd190366760960, 64'd8101555712, - 64'd5013775360, - 64'd365533728, 64'd185296093184, 64'd12149912576, - 64'd4729367040, - 64'd402526848, 64'd178251268096, 64'd15991135232, - 64'd4394157056, - 64'd434266688, 64'd169346187264, 64'd19584544768, - 64'd4012854528, - 64'd460462816, 64'd158714167296, 64'd22892994560, - 64'd3590626816, - 64'd480894272, 64'd146506186752, 64'd25883242496, - 64'd3133030656, - 64'd495411008, 64'd132888772608, 64'd28526272512, - 64'd2645941760, - 64'd503934304, 64'd118041862144, 64'd30797553664, - 64'd2135481216, - 64'd506456576, 64'd102156492800, 64'd32677253120, - 64'd1607940736, - 64'd503040352, 64'd85432393728, 64'd34150387712, - 64'd1069706688, - 64'd493816192, 64'd68075581440, 64'd35206914048, - 64'd527184576, - 64'd478980192, 64'd50295820288, 64'd35841761280, 64'd13275691, - 64'd458790528, 64'd32304191488, 64'd36054810624, 64'd545452224, - 64'd433563520, 64'd14310600704, 64'd35850821632, 64'd1063321216, - 64'd403668896, - 64'd3478606336, 64'd35239272448, 64'd1561123456, - 64'd369524608, - 64'd20862973952, 64'd34234189824, 64'd2033426688, - 64'd331591296, - 64'd37650149376, 64'd32853913600, 64'd2475182848, - 64'd290366144, - 64'd53657956352, 64'd31120795648, 64'd2881780480, - 64'd246376544, - 64'd68716351488, 64'd29060892672, 64'd3249091072, - 64'd200173424, - 64'd82669150208, 64'd26703589376, 64'd3573507840, - 64'd152324528, - 64'd95375622144, 64'd24081211392, 64'd3851980032, - 64'd103407576, - 64'd106711851008, 64'd21228597248, 64'd4082038528, - 64'd54003312, - 64'd116571865088, 64'd18182653952, 64'd4261814272, - 64'd4688806, - 64'd124868567040, 64'd14981902336, 64'd4390051328, 64'd43969216, - 64'd131534446592, 64'd11665993728, 64'd4466109440, 64'd91420760, - 64'd136521965568, 64'd8275239936, 64'd4489962496, 64'd137138640, - 64'd139803836416, 64'd4850135552, 64'd4462188544, 64'd180624272, - 64'd141372964864, 64'd1430882688, 64'd4383951872, 64'd221412864, - 64'd141242171392, - 64'd1943064960, 64'd4256981760, 64'd259078384, - 64'd139443732480, - 64'd5233448448, 64'd4083541248, 64'd293237696, - 64'd136028684288, - 64'd8403623936, 64'd3866393344, 64'd323554464, - 64'd131065856000, - 64'd11418961920, 64'd3608760064, 64'd349742080, - 64'd124640845824, - 64'd14247211008, 64'd3314277632, 64'd371566368, - 64'd116854710272, - 64'd16858833920, 64'd2986947328, 64'd388847200, - 64'd107822514176, - 64'd19227299840, 64'd2631084288, 64'd401459936, - 64'd97671798784, - 64'd21329344512, 64'd2251260672, 64'd409335712, - 64'd86540869632, - 64'd23145181184, 64'd1852249216, 64'd412461504, - 64'd74577018880, - 64'd24658677760, 64'd1438965504, 64'd410879232, - 64'd61934665728, - 64'd25857468416, 64'd1016407424, 64'd404684448, - 64'd48773451776, - 64'd26733047808, 64'd589596736, 64'd394024256, - 64'd35256303616, - 64'd27280797696, 64'd163520480, 64'd379094880, - 64'd21547479040, - 64'd27499972608, - 64'd256926192, 64'd360138432, - 64'd7810651136, - 64'd27393648640, - 64'd666995136, 64'd337439520, 64'd5792974336, - 64'd26968619008, - 64'd1062137472, 64'd311321088, 64'd19106494464, - 64'd26235260928, - 64'd1438052992, 64'd282140192, 64'd31979048960, - 64'd25207339008, - 64'd1790736000, 64'd250283168, 64'd44267466752, - 64'd23901808640, - 64'd2116516096, 64'd216160832, 64'd55837798400, - 64'd22338547712, - 64'd2412095488, 64'd180203184, 64'd66566709248, - 64'd20540094464, - 64'd2674580480, 64'd142854208, 64'd76342730752, - 64'd18531325952, - 64'd2901509120, 64'd104566496, 64'd85067358208, - 64'd16339141632, - 64'd3090871296, 64'd65795828, 64'd92655960064, - 64'd13992113152, - 64'd3241124864, 64'd26995910, 64'd99038543872, - 64'd11520123904, - 64'd3351205888, - 64'd11386859, 64'd104160296960, - 64'd8954007552, - 64'd3420532224, - 64'd48918428, 64'd107981996032, - 64'd6325167616, - 64'd3449003264, - 64'd85181896, 64'd110480179200, - 64'd3665207808, - 64'd3436992256, - 64'd119782032, 64'd111647170560, - 64'd1005561408, - 64'd3385333760, - 64'd152349504, 64'd111490867200, 64'd1622868352, - 64'd3295307008, - 64'd182544688, 64'd110034436096, 64'd4190059008, - 64'd3168613632, - 64'd210061120, 64'd107315757056, 64'd6667201024, - 64'd3007350016, - 64'd234628432, 64'd103386734592, 64'd9027011584, - 64'd2813977088, - 64'd256014944, 64'd98312503296, 64'd11244024832, - 64'd2591285760, - 64'd274029632, 64'd92170379264, 64'd13294855168, - 64'd2342358784, - 64'd288523648, 64'd85048827904, 64'd15158435840, - 64'd2070530560, - 64'd299391392, 64'd77046226944, 64'd16816222208, - 64'd1779343616, - 64'd306570976, 64'd68269547520, 64'd18252363776, - 64'd1472505088, - 64'd310044160, 64'd58832982016, 64'd19453847552, - 64'd1153840384, - 64'd309835904, 64'd48856506368, 64'd20410593280, - 64'd827246976, - 64'd306013216, 64'd38464389120, 64'd21115523072, - 64'd496648352, - 64'd298683904, 64'd27783663616, 64'd21564604416, - 64'd165947968, - 64'd287994368, 64'd16942639104, 64'd21756829696, 64'd161015488, - 64'd274127456, 64'd6069367296, 64'd21694183424, 64'd480511552, - 64'd257299680, - 64'd4709823488, 64'd21381576704, 64'd788959168, - 64'd237758064, - 64'd15271768064, 64'd20826730496, 64'd1082965888, - 64'd215776896, - 64'd25497839616, 64'd20040044544, 64'd1359363712, - 64'd191653968, - 64'd35275247616, 64'd19034429440, 64'd1615242112, - 64'd165706880, - 64'd44498239488, 64'd17825124352, 64'd1847977472, - 64'd138268864, - 64'd53069225984, 64'd16429464576, 64'd2055258368, - 64'd109684824, - 64'd60899762176, 64'd14866663424, 64'd2235107584, - 64'd80307000, - 64'd67911417856, 64'd13157547008, 64'd2385898752, - 64'd50490892, - 64'd74036527104, 64'd11324291072, 64'd2506369792, - 64'd20591002, - 64'd79218802688, 64'd9390139392, 64'd2595631104, 64'd9043209, - 64'd83413778432, 64'd7379118592, 64'd2653169920, 64'd38071296, - 64'd86589120512, 64'd5315746304, 64'd2678849792, 64'd66165620, - 64'd88724840448, 64'd3224739072, 64'd2672905216, 64'd93014920, - 64'd89813286912, 64'd1130721792, 64'd2635934208, 64'd118327656, - 64'd89859039232, - 64'd942053824, 64'd2568883456, 64'd141835040, - 64'd88878645248, - 64'd2969985280, 64'd2473032960, 64'd163293760, - 64'd86900252672, - 64'd4930381312, 64'd2349974784, 64'd182488384, - 64'd83963068416, - 64'd6801708544, 64'd2201590016, 64'd199233408, - 64'd80116711424, - 64'd8563822592, 64'd2030020992, 64'd213374832, - 64'd75420508160, - 64'd10198177792, 64'd1837643904, 64'd224791472, - 64'd69942599680, - 64'd11688014848, 64'd1627035520, 64'd233395808, - 64'd63759036416, - 64'd13018524672, 64'd1400941312, 64'd239134400, - 64'd56952745984, - 64'd14176988160, 64'd1162240128, 64'd241988000, - 64'd49612476416, - 64'd15152887808, 64'd913908864, 64'd241971088, - 64'd41831669760, - 64'd15937992704, 64'd658986304, 64'd239131280, - 64'd33707284480, - 64'd16526415872, 64'd400536864, 64'd233548080, - 64'd25338644480, - 64'd16914642944, 64'd141614768, 64'd225331520, - 64'd16826230784, - 64'd17101535232, - 64'd114771248, 64'd214620368, - 64'd8270504960, - 64'd17088299008, - 64'd365691968, 64'd201579968, 64'd229250672, - 64'd16878435328, - 64'd608330368, 64'd186399968, 64'd8576060928, - 64'd16477662208, - 64'd840012160, 64'd169291648, 64'd16676343808, - 64'd15893807104, - 64'd1058234624, 64'd150485136, 64'd24440932352, - 64'd15136688128, - 64'd1260692480, 64'd130226448, 64'd31786033152, - 64'd14217958400, - 64'd1445301760, 64'd108774312, 64'd38634110976, - 64'd13150946304, - 64'd1610219392, 64'd86397032, 64'd44914671616, - 64'd11950475264, - 64'd1753861248, 64'd63369172, 64'd50564964352, - 64'd10632657920, - 64'd1874915968, 64'd39968276, 64'd55530573824, - 64'd9214700544, - 64'd1972355584, 64'd16471616, 64'd59765919744, - 64'd7714673664, - 64'd2045442560, - 64'd6847026, 64'd63234625536, - 64'd6151298560, - 64'd2093733376, - 64'd29720462, 64'd65909788672, - 64'd4543711744, - 64'd2117079296, - 64'd51891092, 64'd67774132224, - 64'd2911243008, - 64'd2115622528, - 64'd73113720, 64'd68820041728, - 64'd1273183616, - 64'd2089790208, - 64'd93158192, 64'd69049499648, 64'd351433280, - 64'd2040284416, - 64'd111811808, 64'd68473896960, 64'd1944049536, - 64'd1968069376, - 64'd128881496, 64'd67113725952, 64'd3486789120, - 64'd1874356352, - 64'd144195728, 64'd64998219776, 64'd4962652672, - 64'd1760584960, - 64'd157606112, 64'd62164844544, 64'd6355700736, - 64'd1628403200, - 64'd168988784, 64'd58658750464, 64'd7651218944, - 64'd1479644416, - 64'd178245392, 64'd54532087808, 64'd8835868672, - 64'd1316303360, - 64'd185303792, 64'd49843318784, 64'd9897820160, - 64'd1140510208, - 64'd190118496, 64'd44656418816, 64'd10826858496, - 64'd954503680, - 64'd192670752, 64'd39040032768, 64'd11614480384, - 64'd760603392, - 64'd192968256, 64'd33066635264, 64'd12253963264, - 64'd561181504, - 64'd191044672, 64'd26811590656, 64'd12740410368, - 64'd358634592, - 64'd186958800, 64'd20352258048, 64'd13070778368, - 64'd155355344, - 64'd180793488, 64'd13767048192, 64'd13243881472, 64'd46295076, - 64'd172654240, 64'd7134508032, 64'd13260374016, 64'd244013680, - 64'd162667648, 64'd532402080, 64'd13122712576, 64'd435581472, - 64'd150979568, - 64'd5963171840, 64'd12835095552, 64'd618887680, - 64'd137753088, - 64'd12278635520, 64'd12403388416, 64'd791952384, - 64'd123166384, - 64'd18343737344, 64'd11835023360, 64'd952947136, - 64'd107410400, - 64'd24092315648, 64'd11138892800, 64'd1100213760, - 64'd90686408, - 64'd29462990848, 64'd10325217280, 64'd1232280576, - 64'd73203528, - 64'd34399793152, 64'd9405405184, 64'd1347876480, - 64'd55176152, - 64'd38852730880, 64'd8391904768, 64'd1445942016, - 64'd36821416, - 64'd42778251264, 64'd7298036736, 64'd1525638272, - 64'd18356602, - 64'd46139658240, 64'd6137830912, 64'd1586352896, 64'd3364, - 64'd48907403264, 64'd4925849088, 64'd1627703296, 64'd18048354, - 64'd51059314688, 64'd3677007104, 64'd1649537408, 64'd35575396, - 64'd52580737024, 64'd2406398464, 64'd1651931392, 64'd52390896, - 64'd53464559616, 64'd1129114624, 64'd1635185152, 64'd68312728, - 64'd53711183872, - 64'd139928944, 64'd1599814784, 64'd83172152, - 64'd53328396288, - 64'd1386162304, 64'd1546543488, 64'd96815528, - 64'd52331134976, - 64'd2595524096, 64'd1476289152, 64'd109105848, - 64'd50741219328, - 64'd3754616064, 64'd1390150784, 64'd119924056, - 64'd48586973184, - 64'd4850846208, 64'd1289392896, 64'd129170104, - 64'd45902774272, - 64'd5872562688, 64'd1175427840, 64'd136763808, - 64'd42728583168, - 64'd6809170432, 64'd1049796992, 64'd142645424, - 64'd39109353472, - 64'd7651239424, 64'd914150976, 64'd146776032, - 64'd35094458368, - 64'd8390590464, 64'd770228544, 64'd149137584, - 64'd30737025024, - 64'd9020372992, 64'd619834944, 64'd149732832, - 64'd26093264896, - 64'd9535118336, 64'd464820192, 64'd148584864, - 64'd21221765120, - 64'd9930782720, 64'd307056544, 64'd145736576, - 64'd16182777856, - 64'd10204768256, 64'd148416656, 64'd141249808, - 64'd11037487104, - 64'd10355931136, - 64'd9248055, 64'd135204288, - 64'd5847291392, - 64'd10384567296, - 64'd164128624, 64'd127696448, - 64'd673083584, - 64'd10292387840, - 64'd314478656, 64'd118838032, 64'd4425443328, - 64'd10082473984, - 64'd458633504, 64'd108754496, 64'd9390467072, - 64'd9759219712, - 64'd595028224, 64'd97583376, 64'd14166675456, - 64'd9328256000, - 64'd722214016, 64'd85472480, 64'd18701864960, - 64'd8796367872, - 64'd838872960, 64'd72578000, 64'd22947489792, - 64'd8171397632, - 64'd943831040, 64'd59062548, 64'd26859171840, - 64'd7462130688, - 64'd1036069504, 64'd45093212, 64'd30397132800, - 64'd6678184448, - 64'd1114734080, 64'd30839494, 64'd33526589440, - 64'd5829879808, - 64'd1179141760, 64'd16471352, 64'd36218060800, - 64'd4928109056, - 64'd1228786048, 64'd2157196, 64'd38447636480, - 64'd3984203008, - 64'd1263340160, - 64'd11938022, 64'd40197140480, - 64'd3009790464, - 64'd1282657280, - 64'd25654662, 64'd41454268416, - 64'd2016659712, - 64'd1286769408, - 64'd38840152, 64'd42212614144, - 64'd1016618176, - 64'd1275884288, - 64'd51350640, 64'd42471653376, - 64'd21356334, - 64'd1250379776, - 64'd63052516, 64'd42236645376, 64'd957685888, - 64'd1210796416, - 64'd73823768, 64'd41518489600, 64'd1909447296, - 64'd1157828864, - 64'd83555224, 64'd40333484032, 64'd2823367424, - 64'd1092315392, - 64'd92151592, 64'd38703067136, 64'd3689500160, - 64'd1015224960, - 64'd99532312, 64'd36653469696, 64'd4498618368, - 64'd927644736, - 64'd105632264, 64'd34215340032, 64'd5242309120, - 64'd830765056, - 64'd110402272, 64'd31423309824, 64'd5913057792, - 64'd725863872, - 64'd113809368, 64'd28315527168, 64'd6504319488, - 64'd614290688, - 64'd115836928, 64'd24933158912, 64'd7010576896, - 64'd497449664, - 64'd116484592, 64'd21319860224, 64'd7427391488, - 64'd376782464, - 64'd115767992, 64'd17521235968, 64'd7751432704, - 64'd253750912, - 64'd113718288, 64'd13584269312, 64'd7980498432, - 64'd129819680, - 64'd110381560, 64'd9556759552, 64'd8113524224, - 64'd6439408, - 64'd105818040, 64'd5486758400, 64'd8150574080, 64'd114969968, - 64'd100101136, 64'd1422006400, 64'd8092821504, 64'd233035072, - 64'd93316416, - 64'd2590614528, 64'd7942518272, 64'd346444256, - 64'd85560352, - 64'd6505608704, 64'd7702948864, 64'd453961664, - 64'd76939064, - 64'd10279368704, 64'd7378376192, 64'd554440448, - 64'd67566928, - 64'd13870651392, 64'd6973975552, 64'd646834304, - 64'd57565096, - 64'd17241012224, 64'd6495759872, 64'd730208128, - 64'd47059976, - 64'd20355205120, 64'd5950494720, 64'd803746816, - 64'd36181704, - 64'd23181537280, 64'd5345609216, 64'd866762944, - 64'd25062552, - 64'd25692176384, 64'd4689098240, 64'd918702144, - 64'd13835381, - 64'd27863408640, 64'd3989420544, 64'd959147840, - 64'd2632072, - 64'd29675841536, 64'd3255392000, 64'd987823232, 64'd8417969, - 64'd31114557440, 64'd2496078848, 64'd1004592512, 64'd19189274, - 64'd32169211904, 64'd1720688896, 64'd1009460096, 64'd29561700, - 64'd32834078720, 64'd938460864, 64'd1002568000, 64'd39421732, - 64'd33108035584, 64'd158558640, 64'd984192000, 64'd48663680, - 64'd32994498560, - 64'd610034432, 64'd954736192, 64'd57190776};
endpackage
`endif
