`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam N = 4;
	localparam M = 4;
	localparam COEFF_BIAS = 48;
	localparam logic signed[63:0] Lfr[0:3] = {64'd195460265159054, 64'd195460265159054, 64'd218844508241820, 64'd218844508241820};
	localparam logic signed[63:0] Lfi[0:3] = {64'd149205040781794, - 64'd149205040781794, 64'd55594741694325, - 64'd55594741694325};
	localparam logic signed[63:0] Lbr[0:3] = {64'd195460265159054, 64'd195460265159054, 64'd218844508241820, 64'd218844508241820};
	localparam logic signed[63:0] Lbi[0:3] = {64'd149205040781794, - 64'd149205040781794, 64'd55594741694325, - 64'd55594741694325};
	localparam logic signed[63:0] Wfr[0:3] = {64'd71535633211341, 64'd71535633211341, - 64'd3081067831406, - 64'd3081067831406};
	localparam logic signed[63:0] Wfi[0:3] = {- 64'd5570152617347, 64'd5570152617347, - 64'd70391449602042, 64'd70391449602042};
	localparam logic signed[63:0] Wbr[0:3] = {- 64'd71535633211341, - 64'd71535633211341, - 64'd3081067831406, - 64'd3081067831406};
	localparam logic signed[63:0] Wbi[0:3] = {64'd5570152617347, - 64'd5570152617347, - 64'd70391449602042, 64'd70391449602042};
	localparam logic signed[63:0] Ffr[0:3][0:79] = '{
		'{64'd50280979506466, - 64'd26041871146154, - 64'd71274850837395, 64'd17105110276254, 64'd26712956754846, - 64'd58936791093295, - 64'd35047768915953, 64'd32634560356965, - 64'd1274675068037, - 64'd61977976186890, 64'd5721551544869, 64'd32269210390142, - 64'd22157608921632, - 64'd41096289269038, 64'd34694679504023, 64'd19909740103447, - 64'd29800292716169, - 64'd9774173235828, 64'd43818284384230, 64'd3023387614943, - 64'd24476835867944, 64'd17789997033223, 64'd34377144698366, - 64'd10996127468387, - 64'd11250577015756, 64'd32166898588527, 64'd14301892094399, - 64'd17579184183102, 64'd3055573792986, 64'd31097003365379, - 64'd6373726221947, - 64'd16022241598172, 64'd12830098470356, 64'd18638664350887, - 64'd19767204656841, - 64'd8835732306963, 64'd15486798118930, 64'd2152708414137, - 64'd22588839565349, - 64'd43158963025, 64'd11716590796995, - 64'd11235267920090, - 64'd16285716949220, 64'd6683482216735, 64'd4452827920973, - 64'd17246807758587, - 64'd5378290143028, 64'd9315150901538, - 64'd2757875844882, - 64'd15378115906652, 64'd4959720137262, 64'd7836321690034, - 64'd7228611267010, - 64'd8194821426253, 64'd10992907748449, 64'd3773994139697, - 64'd7934494637323, 64'd355360347424, 64'd11482012181579, - 64'd739241943898, - 64'd5502784643442, 64'd6747814694640, 64'd7556771327057, - 64'd3906989233184, - 64'd1586826449136, 64'd9100348129577, 64'd1732000068070, - 64'd4861950078305, 64'd1995889948808, 64'd7488898945287, - 64'd3361869371933, - 64'd3770605356808, 64'd3983013733911, 64'd3455420729858, - 64'd5990921551420, - 64'd1526089246329, 64'd4008462507221, - 64'd916533129936, - 64'd5754588325240, 64'd758245910413},
		'{64'd50280979506466, - 64'd26041871146154, - 64'd71274850837395, 64'd17105110276254, 64'd26712956754846, - 64'd58936791093295, - 64'd35047768915953, 64'd32634560356965, - 64'd1274675068037, - 64'd61977976186890, 64'd5721551544869, 64'd32269210390142, - 64'd22157608921632, - 64'd41096289269038, 64'd34694679504023, 64'd19909740103447, - 64'd29800292716169, - 64'd9774173235828, 64'd43818284384230, 64'd3023387614943, - 64'd24476835867944, 64'd17789997033223, 64'd34377144698366, - 64'd10996127468387, - 64'd11250577015756, 64'd32166898588527, 64'd14301892094399, - 64'd17579184183102, 64'd3055573792986, 64'd31097003365379, - 64'd6373726221947, - 64'd16022241598172, 64'd12830098470356, 64'd18638664350887, - 64'd19767204656841, - 64'd8835732306963, 64'd15486798118930, 64'd2152708414137, - 64'd22588839565349, - 64'd43158963025, 64'd11716590796995, - 64'd11235267920090, - 64'd16285716949220, 64'd6683482216735, 64'd4452827920973, - 64'd17246807758587, - 64'd5378290143028, 64'd9315150901538, - 64'd2757875844882, - 64'd15378115906652, 64'd4959720137262, 64'd7836321690034, - 64'd7228611267010, - 64'd8194821426253, 64'd10992907748449, 64'd3773994139697, - 64'd7934494637323, 64'd355360347424, 64'd11482012181579, - 64'd739241943898, - 64'd5502784643442, 64'd6747814694640, 64'd7556771327057, - 64'd3906989233184, - 64'd1586826449136, 64'd9100348129577, 64'd1732000068070, - 64'd4861950078305, 64'd1995889948808, 64'd7488898945287, - 64'd3361869371933, - 64'd3770605356808, 64'd3983013733911, 64'd3455420729858, - 64'd5990921551420, - 64'd1526089246329, 64'd4008462507221, - 64'd916533129936, - 64'd5754588325240, 64'd758245910413},
		'{- 64'd11487437080834, - 64'd47131574021965, - 64'd393791824171, - 64'd69410655546100, - 64'd25067534052799, - 64'd33970843015857, - 64'd9880246262373, - 64'd51571859639094, - 64'd31587388625152, - 64'd22494720173892, - 64'd15110215557093, - 64'd35527321679727, - 64'd32986800495394, - 64'd13118527688908, - 64'd17138154939844, - 64'd22057674596806, - 64'd30967306231497, - 64'd5923639544567, - 64'd16926057972688, - 64'd11437327597160, - 64'd26926497355389, - 64'd769329185019, - 64'd15291262131942, - 64'd3590641589677, - 64'd21942659220809, 64'd2615595438176, - 64'd12885666548256, 64'd1776584594975, - 64'd16793151339178, 64'd4562275356497, - 64'd10197003281649, 64'd5073154886266, - 64'd11992873441878, 64'd5411116139979, - 64'd7564187615261, 64'd6745432921861, - 64'd7842251756373, 64'd5478352113918, - 64'd5200369441332, 64'd7224439661996, - 64'd4477103794630, 64'd5036669936686, - 64'd3218899805939, 64'd6893168604395, - 64'd1915297895408, 64'd4306594661297, - 64'd1658874789301, 64'd6069804407600, - 64'd97219829399, 64'd3455564019637, - 64'd508146231406, 64'd5002660935327, 64'd1081327921369, 64'd2602032059218, 64'd277334570179, 64'd3873108892229, 64'd1744008768652, 64'd1822445934134, 64'd758245234275, 64'd2803385642161, 64'd2016065717516, 64'd1159453992167, 64'd1000592925925, 64'd1866855401359, 64'd2012671621041, 64'd630179619198, 64'd1067971382313, 64'd1098938017507, 64'd1832323933842, 64'd233804990339, 64'd1016791911511, 64'd507500561226, 64'd1554070326828, - 64'd41960577938, 64'd893850313143, 64'd81983361463, 64'd1237445070286, - 64'd215702624716, 64'd735612354203, - 64'd199096195571},
		'{- 64'd11487437080834, - 64'd47131574021965, - 64'd393791824171, - 64'd69410655546099, - 64'd25067534052799, - 64'd33970843015857, - 64'd9880246262373, - 64'd51571859639094, - 64'd31587388625152, - 64'd22494720173892, - 64'd15110215557093, - 64'd35527321679727, - 64'd32986800495394, - 64'd13118527688908, - 64'd17138154939844, - 64'd22057674596806, - 64'd30967306231497, - 64'd5923639544567, - 64'd16926057972688, - 64'd11437327597160, - 64'd26926497355389, - 64'd769329185019, - 64'd15291262131942, - 64'd3590641589677, - 64'd21942659220809, 64'd2615595438176, - 64'd12885666548256, 64'd1776584594975, - 64'd16793151339178, 64'd4562275356497, - 64'd10197003281649, 64'd5073154886266, - 64'd11992873441878, 64'd5411116139979, - 64'd7564187615261, 64'd6745432921861, - 64'd7842251756373, 64'd5478352113918, - 64'd5200369441332, 64'd7224439661996, - 64'd4477103794630, 64'd5036669936686, - 64'd3218899805939, 64'd6893168604395, - 64'd1915297895408, 64'd4306594661297, - 64'd1658874789301, 64'd6069804407600, - 64'd97219829399, 64'd3455564019637, - 64'd508146231406, 64'd5002660935327, 64'd1081327921369, 64'd2602032059218, 64'd277334570179, 64'd3873108892229, 64'd1744008768652, 64'd1822445934134, 64'd758245234275, 64'd2803385642161, 64'd2016065717516, 64'd1159453992167, 64'd1000592925925, 64'd1866855401359, 64'd2012671621041, 64'd630179619198, 64'd1067971382313, 64'd1098938017507, 64'd1832323933842, 64'd233804990339, 64'd1016791911511, 64'd507500561226, 64'd1554070326828, - 64'd41960577938, 64'd893850313143, 64'd81983361463, 64'd1237445070286, - 64'd215702624716, 64'd735612354203, - 64'd199096195571}};
	localparam logic signed[63:0] Ffi[0:3][0:79] = '{
		'{64'd15474709797000, 64'd77068983733182, - 64'd27253310499194, - 64'd39157140373105, 64'd37398942531268, 64'd39713461140531, - 64'd56706661846364, - 64'd18124155914208, 64'd40130441284130, - 64'd3663781007330, - 64'd57956139269744, 64'd4713344694742, 64'd27191471292682, - 64'd35397640629197, - 64'd37212679223131, 64'd20378367281913, 64'd7136780930328, - 64'd46365065528260, - 64'd7449966254295, 64'd24704841395792, - 64'd10840739140155, - 64'd37377688210436, 64'd18053954878804, 64'd18758042309914, - 64'd20502714337811, - 64'd16525432101113, 64'd30759658231936, 64'd7196995981922, - 64'd20201116453946, 64'd5575622009863, 64'd28941135168089, - 64'd4320725643848, - 64'd12408238227845, 64'd20355778260486, 64'd16718537214477, - 64'd11493488440440, - 64'd1815444394521, 64'd24015379874618, 64'd1131337299565, - 64'd12664913020076, 64'd6948614491547, 64'd17817738271158, - 64'd11188338220350, - 64'd8817575263573, 64'd11035980800127, 64'd6417271119133, - 64'd16402120965637, - 64'd2580251967166, 64'd10023910963590, - 64'd4685990761404, - 64'd14240807335998, 64'd3146037160466, 64'd5498845172864, - 64'd11405693839194, - 64'd7259958794588, 64'd6338552633614, - 64'd13285384645, - 64'd12264211361083, 64'd785731578944, 64'd6402111296263, - 64'd4215164611132, - 64'd8328074050732, 64'd6632040334060, 64'd4053858572058, - 64'd5844002258894, - 64'd2206233757528, 64'd8611098452154, 64'd744029845878, - 64'd4899308465306, 64'd3291897522760, 64'd6897773827885, - 64'd2060571051569, - 64'd2344163229811, 64'd6255677345796, 64'd3007844088157, - 64'd3429623128260, 64'd483506426462, 64'd6175691224810, - 64'd1086994286126, - 64'd3190533186201},
		'{- 64'd15474709797000, - 64'd77068983733182, 64'd27253310499194, 64'd39157140373105, - 64'd37398942531268, - 64'd39713461140531, 64'd56706661846364, 64'd18124155914208, - 64'd40130441284130, 64'd3663781007330, 64'd57956139269744, - 64'd4713344694742, - 64'd27191471292682, 64'd35397640629197, 64'd37212679223131, - 64'd20378367281913, - 64'd7136780930328, 64'd46365065528260, 64'd7449966254295, - 64'd24704841395792, 64'd10840739140155, 64'd37377688210436, - 64'd18053954878804, - 64'd18758042309914, 64'd20502714337811, 64'd16525432101113, - 64'd30759658231936, - 64'd7196995981922, 64'd20201116453946, - 64'd5575622009863, - 64'd28941135168089, 64'd4320725643848, 64'd12408238227845, - 64'd20355778260486, - 64'd16718537214477, 64'd11493488440440, 64'd1815444394521, - 64'd24015379874618, - 64'd1131337299565, 64'd12664913020076, - 64'd6948614491547, - 64'd17817738271158, 64'd11188338220350, 64'd8817575263573, - 64'd11035980800127, - 64'd6417271119133, 64'd16402120965637, 64'd2580251967166, - 64'd10023910963590, 64'd4685990761404, 64'd14240807335998, - 64'd3146037160466, - 64'd5498845172864, 64'd11405693839194, 64'd7259958794588, - 64'd6338552633614, 64'd13285384645, 64'd12264211361083, - 64'd785731578944, - 64'd6402111296263, 64'd4215164611132, 64'd8328074050732, - 64'd6632040334060, - 64'd4053858572058, 64'd5844002258894, 64'd2206233757528, - 64'd8611098452154, - 64'd744029845878, 64'd4899308465306, - 64'd3291897522760, - 64'd6897773827885, 64'd2060571051569, 64'd2344163229811, - 64'd6255677345796, - 64'd3007844088157, 64'd3429623128260, - 64'd483506426462, - 64'd6175691224810, 64'd1086994286126, 64'd3190533186201},
		'{64'd81696953819194, - 64'd13536242274637, 64'd48473341657088, - 64'd12122599518399, 64'd61249809086581, - 64'd19833379267571, 64'd37609850746766, - 64'd23134673896180, 64'd42670085310018, - 64'd22129947208747, 64'd27289884318162, - 64'd28173092472186, 64'd26936750163365, - 64'd21648835868395, 64'd18233211501489, - 64'd28921430013904, 64'd14427808957402, - 64'd19422863310231, 64'd10791179177668, - 64'd26842836755599, 64'd5101083521384, - 64'd16271109544683, 64'd5046951228818, - 64'd23129099286592, - 64'd1352260705076, - 64'd12802607415715, 64'd903752775321, - 64'd18691882357108, - 64'd5385314595986, - 64'd9437311275004, - 64'd1842415896726, - 64'd14181889585883, - 64'd7503890612602, - 64'd6436327826692, - 64'd3446495939824, - 64'd10024293988256, - 64'd8202952813680, - 64'd3935431159745, - 64'd4173641932347, - 64'd6461501866625, - 64'd7926669579696, - 64'd1977724388489, - 64'd4272109109379, - 64'd3596850254475, - 64'd7047203834408, - 64'd542860892619, - 64'd3957302114261, - 64'd1435036967988, - 64'd5857438443200, 64'd428535048116, - 64'd3404418260452, 64'd83130830601, - 64'd4573312917564, 64'd1015698568627, - 64'd2747272626408, 64'd1052720109223, - 64'd3342138192880, 64'd1303630462195, - 64'd2081205192683, 64'd1583467590069, - 64'd2254022292516, 64'd1373517400751, - 64'd1468357449861, 64'd1784836053925, - 64'd1354286451401, 64'd1296904931287, - 64'd944006681820, 64'd1756422251492, - 64'd655419518083, 64'd1132801213097, - 64'd523020151360, 64'd1582657699523, - 64'd147677021988, 64'd926923080373, - 64'd205815113033, 64'd1330741058959, 64'd192130162941, 64'd712387440453, 64'd16526762437, 64'd1050833079037},
		'{- 64'd81696953819194, 64'd13536242274637, - 64'd48473341657088, 64'd12122599518399, - 64'd61249809086581, 64'd19833379267571, - 64'd37609850746766, 64'd23134673896180, - 64'd42670085310018, 64'd22129947208747, - 64'd27289884318162, 64'd28173092472186, - 64'd26936750163365, 64'd21648835868395, - 64'd18233211501489, 64'd28921430013904, - 64'd14427808957402, 64'd19422863310231, - 64'd10791179177668, 64'd26842836755598, - 64'd5101083521384, 64'd16271109544683, - 64'd5046951228818, 64'd23129099286592, 64'd1352260705076, 64'd12802607415715, - 64'd903752775321, 64'd18691882357108, 64'd5385314595986, 64'd9437311275004, 64'd1842415896726, 64'd14181889585883, 64'd7503890612602, 64'd6436327826692, 64'd3446495939824, 64'd10024293988256, 64'd8202952813680, 64'd3935431159745, 64'd4173641932347, 64'd6461501866625, 64'd7926669579696, 64'd1977724388489, 64'd4272109109379, 64'd3596850254475, 64'd7047203834408, 64'd542860892619, 64'd3957302114261, 64'd1435036967988, 64'd5857438443200, - 64'd428535048116, 64'd3404418260452, - 64'd83130830601, 64'd4573312917564, - 64'd1015698568627, 64'd2747272626408, - 64'd1052720109223, 64'd3342138192880, - 64'd1303630462195, 64'd2081205192683, - 64'd1583467590069, 64'd2254022292516, - 64'd1373517400751, 64'd1468357449861, - 64'd1784836053925, 64'd1354286451401, - 64'd1296904931287, 64'd944006681820, - 64'd1756422251492, 64'd655419518083, - 64'd1132801213097, 64'd523020151360, - 64'd1582657699523, 64'd147677021988, - 64'd926923080373, 64'd205815113033, - 64'd1330741058959, - 64'd192130162941, - 64'd712387440453, - 64'd16526762437, - 64'd1050833079037}};
	localparam logic signed[63:0] Fbr[0:3][0:79] = '{
		'{- 64'd50280979506466, - 64'd26041871146154, 64'd71274850837395, 64'd17105110276254, - 64'd26712956754846, - 64'd58936791093295, 64'd35047768915953, 64'd32634560356965, 64'd1274675068037, - 64'd61977976186890, - 64'd5721551544869, 64'd32269210390142, 64'd22157608921632, - 64'd41096289269038, - 64'd34694679504023, 64'd19909740103447, 64'd29800292716169, - 64'd9774173235828, - 64'd43818284384230, 64'd3023387614943, 64'd24476835867944, 64'd17789997033223, - 64'd34377144698366, - 64'd10996127468387, 64'd11250577015756, 64'd32166898588527, - 64'd14301892094399, - 64'd17579184183102, - 64'd3055573792986, 64'd31097003365379, 64'd6373726221947, - 64'd16022241598172, - 64'd12830098470356, 64'd18638664350887, 64'd19767204656841, - 64'd8835732306963, - 64'd15486798118930, 64'd2152708414137, 64'd22588839565349, - 64'd43158963025, - 64'd11716590796995, - 64'd11235267920090, 64'd16285716949220, 64'd6683482216735, - 64'd4452827920973, - 64'd17246807758587, 64'd5378290143028, 64'd9315150901538, 64'd2757875844882, - 64'd15378115906652, - 64'd4959720137262, 64'd7836321690034, 64'd7228611267010, - 64'd8194821426253, - 64'd10992907748449, 64'd3773994139697, 64'd7934494637323, 64'd355360347424, - 64'd11482012181579, - 64'd739241943898, 64'd5502784643442, 64'd6747814694640, - 64'd7556771327057, - 64'd3906989233184, 64'd1586826449136, 64'd9100348129577, - 64'd1732000068070, - 64'd4861950078305, - 64'd1995889948808, 64'd7488898945287, 64'd3361869371933, - 64'd3770605356808, - 64'd3983013733911, 64'd3455420729858, 64'd5990921551420, - 64'd1526089246329, - 64'd4008462507221, - 64'd916533129936, 64'd5754588325240, 64'd758245910413},
		'{- 64'd50280979506466, - 64'd26041871146154, 64'd71274850837395, 64'd17105110276254, - 64'd26712956754846, - 64'd58936791093295, 64'd35047768915953, 64'd32634560356965, 64'd1274675068037, - 64'd61977976186890, - 64'd5721551544869, 64'd32269210390142, 64'd22157608921632, - 64'd41096289269038, - 64'd34694679504023, 64'd19909740103447, 64'd29800292716169, - 64'd9774173235828, - 64'd43818284384230, 64'd3023387614943, 64'd24476835867944, 64'd17789997033223, - 64'd34377144698366, - 64'd10996127468387, 64'd11250577015756, 64'd32166898588527, - 64'd14301892094399, - 64'd17579184183102, - 64'd3055573792986, 64'd31097003365379, 64'd6373726221947, - 64'd16022241598172, - 64'd12830098470356, 64'd18638664350887, 64'd19767204656841, - 64'd8835732306963, - 64'd15486798118930, 64'd2152708414137, 64'd22588839565349, - 64'd43158963025, - 64'd11716590796995, - 64'd11235267920090, 64'd16285716949220, 64'd6683482216735, - 64'd4452827920973, - 64'd17246807758587, 64'd5378290143028, 64'd9315150901538, 64'd2757875844882, - 64'd15378115906652, - 64'd4959720137262, 64'd7836321690034, 64'd7228611267010, - 64'd8194821426253, - 64'd10992907748449, 64'd3773994139697, 64'd7934494637323, 64'd355360347424, - 64'd11482012181579, - 64'd739241943898, 64'd5502784643442, 64'd6747814694640, - 64'd7556771327057, - 64'd3906989233184, 64'd1586826449136, 64'd9100348129577, - 64'd1732000068070, - 64'd4861950078305, - 64'd1995889948808, 64'd7488898945287, 64'd3361869371933, - 64'd3770605356808, - 64'd3983013733911, 64'd3455420729858, 64'd5990921551420, - 64'd1526089246329, - 64'd4008462507221, - 64'd916533129936, 64'd5754588325240, 64'd758245910413},
		'{- 64'd11487437080834, 64'd47131574021965, - 64'd393791824171, 64'd69410655546100, - 64'd25067534052799, 64'd33970843015857, - 64'd9880246262373, 64'd51571859639094, - 64'd31587388625152, 64'd22494720173892, - 64'd15110215557093, 64'd35527321679727, - 64'd32986800495394, 64'd13118527688908, - 64'd17138154939844, 64'd22057674596806, - 64'd30967306231497, 64'd5923639544567, - 64'd16926057972688, 64'd11437327597160, - 64'd26926497355389, 64'd769329185019, - 64'd15291262131942, 64'd3590641589677, - 64'd21942659220809, - 64'd2615595438176, - 64'd12885666548256, - 64'd1776584594975, - 64'd16793151339178, - 64'd4562275356497, - 64'd10197003281649, - 64'd5073154886266, - 64'd11992873441878, - 64'd5411116139979, - 64'd7564187615261, - 64'd6745432921861, - 64'd7842251756373, - 64'd5478352113918, - 64'd5200369441332, - 64'd7224439661996, - 64'd4477103794630, - 64'd5036669936686, - 64'd3218899805939, - 64'd6893168604395, - 64'd1915297895408, - 64'd4306594661297, - 64'd1658874789301, - 64'd6069804407600, - 64'd97219829399, - 64'd3455564019637, - 64'd508146231406, - 64'd5002660935327, 64'd1081327921369, - 64'd2602032059218, 64'd277334570179, - 64'd3873108892229, 64'd1744008768652, - 64'd1822445934134, 64'd758245234275, - 64'd2803385642161, 64'd2016065717516, - 64'd1159453992167, 64'd1000592925925, - 64'd1866855401359, 64'd2012671621041, - 64'd630179619198, 64'd1067971382313, - 64'd1098938017507, 64'd1832323933842, - 64'd233804990339, 64'd1016791911511, - 64'd507500561226, 64'd1554070326828, 64'd41960577938, 64'd893850313143, - 64'd81983361463, 64'd1237445070286, 64'd215702624716, 64'd735612354203, 64'd199096195571},
		'{- 64'd11487437080834, 64'd47131574021965, - 64'd393791824171, 64'd69410655546099, - 64'd25067534052799, 64'd33970843015857, - 64'd9880246262373, 64'd51571859639094, - 64'd31587388625152, 64'd22494720173892, - 64'd15110215557093, 64'd35527321679727, - 64'd32986800495394, 64'd13118527688908, - 64'd17138154939844, 64'd22057674596806, - 64'd30967306231497, 64'd5923639544567, - 64'd16926057972688, 64'd11437327597160, - 64'd26926497355389, 64'd769329185019, - 64'd15291262131942, 64'd3590641589677, - 64'd21942659220809, - 64'd2615595438176, - 64'd12885666548256, - 64'd1776584594975, - 64'd16793151339178, - 64'd4562275356497, - 64'd10197003281649, - 64'd5073154886266, - 64'd11992873441878, - 64'd5411116139979, - 64'd7564187615261, - 64'd6745432921861, - 64'd7842251756373, - 64'd5478352113918, - 64'd5200369441332, - 64'd7224439661996, - 64'd4477103794630, - 64'd5036669936686, - 64'd3218899805939, - 64'd6893168604395, - 64'd1915297895408, - 64'd4306594661297, - 64'd1658874789301, - 64'd6069804407600, - 64'd97219829399, - 64'd3455564019637, - 64'd508146231406, - 64'd5002660935327, 64'd1081327921369, - 64'd2602032059218, 64'd277334570179, - 64'd3873108892229, 64'd1744008768652, - 64'd1822445934134, 64'd758245234275, - 64'd2803385642161, 64'd2016065717516, - 64'd1159453992167, 64'd1000592925925, - 64'd1866855401359, 64'd2012671621041, - 64'd630179619198, 64'd1067971382313, - 64'd1098938017507, 64'd1832323933842, - 64'd233804990339, 64'd1016791911511, - 64'd507500561226, 64'd1554070326828, 64'd41960577938, 64'd893850313143, - 64'd81983361463, 64'd1237445070286, 64'd215702624716, 64'd735612354203, 64'd199096195571}};
	localparam logic signed[63:0] Fbi[0:3][0:79] = '{
		'{- 64'd15474709797000, 64'd77068983733182, 64'd27253310499194, - 64'd39157140373105, - 64'd37398942531268, 64'd39713461140531, 64'd56706661846364, - 64'd18124155914208, - 64'd40130441284130, - 64'd3663781007330, 64'd57956139269744, 64'd4713344694742, - 64'd27191471292682, - 64'd35397640629197, 64'd37212679223131, 64'd20378367281913, - 64'd7136780930328, - 64'd46365065528260, 64'd7449966254295, 64'd24704841395792, 64'd10840739140155, - 64'd37377688210436, - 64'd18053954878804, 64'd18758042309914, 64'd20502714337811, - 64'd16525432101113, - 64'd30759658231936, 64'd7196995981922, 64'd20201116453946, 64'd5575622009863, - 64'd28941135168089, - 64'd4320725643848, 64'd12408238227845, 64'd20355778260486, - 64'd16718537214477, - 64'd11493488440440, 64'd1815444394521, 64'd24015379874618, - 64'd1131337299565, - 64'd12664913020076, - 64'd6948614491547, 64'd17817738271158, 64'd11188338220350, - 64'd8817575263573, - 64'd11035980800127, 64'd6417271119133, 64'd16402120965637, - 64'd2580251967166, - 64'd10023910963590, - 64'd4685990761404, 64'd14240807335998, 64'd3146037160466, - 64'd5498845172864, - 64'd11405693839194, 64'd7259958794588, 64'd6338552633614, 64'd13285384645, - 64'd12264211361083, - 64'd785731578944, 64'd6402111296263, 64'd4215164611132, - 64'd8328074050732, - 64'd6632040334060, 64'd4053858572058, 64'd5844002258894, - 64'd2206233757528, - 64'd8611098452154, 64'd744029845878, 64'd4899308465306, 64'd3291897522760, - 64'd6897773827885, - 64'd2060571051569, 64'd2344163229811, 64'd6255677345796, - 64'd3007844088157, - 64'd3429623128260, - 64'd483506426462, 64'd6175691224810, 64'd1086994286126, - 64'd3190533186201},
		'{64'd15474709797000, - 64'd77068983733182, - 64'd27253310499194, 64'd39157140373105, 64'd37398942531268, - 64'd39713461140531, - 64'd56706661846364, 64'd18124155914208, 64'd40130441284130, 64'd3663781007330, - 64'd57956139269744, - 64'd4713344694742, 64'd27191471292682, 64'd35397640629197, - 64'd37212679223131, - 64'd20378367281913, 64'd7136780930328, 64'd46365065528260, - 64'd7449966254295, - 64'd24704841395792, - 64'd10840739140155, 64'd37377688210436, 64'd18053954878804, - 64'd18758042309914, - 64'd20502714337811, 64'd16525432101113, 64'd30759658231936, - 64'd7196995981922, - 64'd20201116453946, - 64'd5575622009863, 64'd28941135168089, 64'd4320725643848, - 64'd12408238227845, - 64'd20355778260486, 64'd16718537214477, 64'd11493488440440, - 64'd1815444394521, - 64'd24015379874618, 64'd1131337299565, 64'd12664913020076, 64'd6948614491547, - 64'd17817738271158, - 64'd11188338220350, 64'd8817575263573, 64'd11035980800127, - 64'd6417271119133, - 64'd16402120965637, 64'd2580251967166, 64'd10023910963590, 64'd4685990761404, - 64'd14240807335998, - 64'd3146037160466, 64'd5498845172864, 64'd11405693839194, - 64'd7259958794588, - 64'd6338552633614, - 64'd13285384645, 64'd12264211361083, 64'd785731578944, - 64'd6402111296263, - 64'd4215164611132, 64'd8328074050732, 64'd6632040334060, - 64'd4053858572058, - 64'd5844002258894, 64'd2206233757528, 64'd8611098452154, - 64'd744029845878, - 64'd4899308465306, - 64'd3291897522760, 64'd6897773827885, 64'd2060571051569, - 64'd2344163229811, - 64'd6255677345796, 64'd3007844088157, 64'd3429623128260, 64'd483506426462, - 64'd6175691224810, - 64'd1086994286126, 64'd3190533186201},
		'{64'd81696953819194, 64'd13536242274637, 64'd48473341657088, 64'd12122599518399, 64'd61249809086581, 64'd19833379267571, 64'd37609850746766, 64'd23134673896180, 64'd42670085310018, 64'd22129947208747, 64'd27289884318162, 64'd28173092472186, 64'd26936750163365, 64'd21648835868395, 64'd18233211501489, 64'd28921430013904, 64'd14427808957402, 64'd19422863310231, 64'd10791179177668, 64'd26842836755599, 64'd5101083521384, 64'd16271109544683, 64'd5046951228818, 64'd23129099286592, - 64'd1352260705076, 64'd12802607415715, 64'd903752775321, 64'd18691882357108, - 64'd5385314595986, 64'd9437311275004, - 64'd1842415896726, 64'd14181889585883, - 64'd7503890612602, 64'd6436327826692, - 64'd3446495939824, 64'd10024293988256, - 64'd8202952813680, 64'd3935431159745, - 64'd4173641932347, 64'd6461501866625, - 64'd7926669579696, 64'd1977724388489, - 64'd4272109109379, 64'd3596850254475, - 64'd7047203834408, 64'd542860892619, - 64'd3957302114261, 64'd1435036967988, - 64'd5857438443200, - 64'd428535048116, - 64'd3404418260452, - 64'd83130830601, - 64'd4573312917564, - 64'd1015698568627, - 64'd2747272626408, - 64'd1052720109223, - 64'd3342138192880, - 64'd1303630462195, - 64'd2081205192683, - 64'd1583467590069, - 64'd2254022292516, - 64'd1373517400751, - 64'd1468357449861, - 64'd1784836053925, - 64'd1354286451401, - 64'd1296904931287, - 64'd944006681820, - 64'd1756422251492, - 64'd655419518083, - 64'd1132801213097, - 64'd523020151360, - 64'd1582657699523, - 64'd147677021988, - 64'd926923080373, - 64'd205815113033, - 64'd1330741058959, 64'd192130162941, - 64'd712387440453, 64'd16526762437, - 64'd1050833079037},
		'{- 64'd81696953819194, - 64'd13536242274637, - 64'd48473341657088, - 64'd12122599518399, - 64'd61249809086581, - 64'd19833379267571, - 64'd37609850746766, - 64'd23134673896180, - 64'd42670085310018, - 64'd22129947208747, - 64'd27289884318162, - 64'd28173092472186, - 64'd26936750163365, - 64'd21648835868395, - 64'd18233211501489, - 64'd28921430013904, - 64'd14427808957402, - 64'd19422863310231, - 64'd10791179177668, - 64'd26842836755598, - 64'd5101083521384, - 64'd16271109544683, - 64'd5046951228818, - 64'd23129099286592, 64'd1352260705076, - 64'd12802607415715, - 64'd903752775321, - 64'd18691882357108, 64'd5385314595986, - 64'd9437311275004, 64'd1842415896726, - 64'd14181889585883, 64'd7503890612602, - 64'd6436327826692, 64'd3446495939824, - 64'd10024293988256, 64'd8202952813680, - 64'd3935431159745, 64'd4173641932347, - 64'd6461501866625, 64'd7926669579696, - 64'd1977724388489, 64'd4272109109379, - 64'd3596850254475, 64'd7047203834408, - 64'd542860892619, 64'd3957302114261, - 64'd1435036967988, 64'd5857438443200, 64'd428535048116, 64'd3404418260452, 64'd83130830601, 64'd4573312917564, 64'd1015698568627, 64'd2747272626408, 64'd1052720109223, 64'd3342138192880, 64'd1303630462195, 64'd2081205192683, 64'd1583467590069, 64'd2254022292516, 64'd1373517400751, 64'd1468357449861, 64'd1784836053925, 64'd1354286451401, 64'd1296904931287, 64'd944006681820, 64'd1756422251492, 64'd655419518083, 64'd1132801213097, 64'd523020151360, 64'd1582657699523, 64'd147677021988, 64'd926923080373, 64'd205815113033, 64'd1330741058959, - 64'd192130162941, 64'd712387440453, - 64'd16526762437, 64'd1050833079037}};
	localparam logic signed[63:0] hf[0:1199] = {64'd67282986336256, - 64'd15925081276416, - 64'd13053910319104, 64'd2600907833344, 64'd46241719255040, - 64'd37561451937792, - 64'd1031533821952, 64'd5428495253504, 64'd22973836689408, - 64'd42223953510400, 64'd14594550530048, 64'd3275386781696, 64'd4008551907328, - 64'd32830579015680, 64'd25656928763904, - 64'd3055999516672, - 64'd6970588266496, - 64'd16388061134848, 64'd27745474052096, - 64'd10660821860352, - 64'd9729572077568, - 64'd558183612416, 64'd21047197827072, - 64'd16336497410048, - 64'd6726005817344, 64'd9235473629184, 64'd9221060952064, - 64'd18038350938112, - 64'd1572290035712, 64'd11206951698432, - 64'd2792537194496, - 64'd15519267684352, 64'd2539725258752, 64'd6941853089792, - 64'd10944011829248, - 64'd10107455799296, 64'd3868836757504, - 64'd43593134080, - 64'd13410579251200, - 64'd3913146171392, 64'd2363855470592, - 64'd6105038061568, - 64'd10786977087488, 64'd1098257989632, - 64'd782689632256, - 64'd8878215397376, - 64'd5325878984704, 64'd3782055559168, - 64'd3932610363392, - 64'd7863339057152, 64'd265721282560, 64'd4039707721728, - 64'd5767671840768, - 64'd4165725585408, 64'd3920110813184, 64'd2610896044032, - 64'd5743348547584, 64'd307357745152, 64'd4809766207488, 64'd608251281408, - 64'd4135357513728, 64'd3761841111040, 64'd3347204800512, - 64'd973607337984, - 64'd1759289540608, 64'd5173173813248, 64'd725637267456, - 64'd1587403030528, 64'd452657709056, 64'd4498294571008, - 64'd1719660838912, - 64'd1217645772800, 64'd1823868452864, 64'd2468478976000, - 64'd3048596832256, - 64'd247646093312, 64'd2125608386560, 64'd139588567040, - 64'd2975866552320, 64'd789078605824, 64'd1558683582464, - 64'd1574487588864, - 64'd1822248665088, 64'd1452403195904, 64'd580105928704, - 64'd2206403395584, - 64'd249477169152, 64'd1544294105088, - 64'd324482531328, - 64'd1802040639488, 64'd1070292205568, 64'd1129679159296, - 64'd825176489984, - 64'd780396658688, 64'd1710814658560, 64'd452293754880, - 64'd830565056512, 64'd312181686272, 64'd1595238514688, - 64'd197752094720, - 64'd462174879744, 64'd1036644909056, 64'd944033038336, - 64'd603327168512, 64'd44093468672, 64'd1199774105600, 64'd123612667904, - 64'd684659245056, 64'd455350353920, 64'd867670949888, - 64'd524179013632, - 64'd497407426560, 64'd629578399744, 64'd278893756416, - 64'd803341008896, - 64'd180656930816, 64'd548160176128, - 64'd286385700864, - 64'd701962387456, 64'd113976459264, 64'd294101155840, - 64'd621751107584, - 64'd352735592448, 64'd281209077760, - 64'd2937806080, - 64'd654878048256, 64'd51129118720, 64'd289786101760, - 64'd226267906048, - 64'd443271741440, 64'd342598811648, 64'd176047620096, - 64'd312955174912, - 64'd122301136896, 64'd437094350848, 64'd13857614848, - 64'd264891580416, 64'd163707863040, 64'd344519704576, - 64'd122259980288, - 64'd132998979584, 64'd317496164352, 64'd143046770688, - 64'd185387843584, 64'd13189578752, 64'd314071711744, - 64'd66452946944, - 64'd167360462848, 64'd115740844032, 64'd192934281216, - 64'd203674533888, - 64'd92692570112, 64'd147073630208, 64'd28029116416, - 64'd234183180288, - 64'd1661353472, 64'd112948879360, - 64'd108060467200, - 64'd171532304384, 64'd68537696256, 64'd42308988928, - 64'd170921951232, - 64'd60893442048, 64'd97036427264, - 64'd29120120832, - 64'd154225328128, 64'd45294145536, 64'd83297353728, - 64'd73854386176, - 64'd83033202688, 64'd108645400576, 64'd42557046784, - 64'd81010794496, 64'd3052362496, 64'd115854442496, - 64'd3562243584, - 64'd56455655424, 64'd68188557312, 64'd77730291712, - 64'd36616466432, - 64'd16636317696, 64'd92843220992, 64'd19440162816, - 64'd47458037760, 64'd20094365696, 64'd77261340672, - 64'd32307419136, - 64'd37433786368, 64'd40815644672, 64'd36701044736, - 64'd59619008512, - 64'd15378306048, 64'd41605963776, - 64'd7827344896, - 64'd58019115008, 64'd7477295104, 64'd26895316992, - 64'd38786220032, - 64'd34939965440, 64'd22283012096, 64'd5842346496, - 64'd47853600768, - 64'd4111832064, 64'd25320962048, - 64'd12203354112, - 64'd36857671680, 64'd21074898944, 64'd18181029888, - 64'd21238448128, - 64'd14691079168, 64'd32507189248, 64'd5906238976, - 64'd20055070720, 64'd7688411648, 64'd29140660224, - 64'd5716253184, - 64'd11553614848, 64'd21846499328, 64'd15719245824, - 64'd12501473280, - 64'd681912448, 64'd24429867008, - 64'd369907456, - 64'd13057359872, 64'd7902852096, 64'd17216260096, - 64'd12487081984, - 64'd8647524352, 64'd11508850688, 64'd5232218624, - 64'd17048470528, - 64'd2091785984, 64'd9951410176, - 64'd5899296256, - 64'd14144353280, 64'd3656101120, 64'd5027585536, - 64'd12206102528, - 64'd6635649536, 64'd6644591616, - 64'd626875840, - 64'd12463518720, 64'd1572722304, 64'd6416714240, - 64'd4723875840, - 64'd8002545664, 64'd7240418816, 64'd3826697984, - 64'd6098137600, - 64'd1606498944, 64'd8846891008, 64'd409438048, - 64'd4878330880, 64'd3874911744, 64'd6752942592, - 64'd2355343360, - 64'd2133099008, 64'd6608261632, 64'd2619789312, - 64'd3583894528, 64'd751143296, 64'd6222286336, - 64'd1521067904, - 64'd3177977344, 64'd2664177920, 64'd3600797952, - 64'd4116261888, - 64'd1675420032, 64'd3122017536, 64'd254774480, - 64'd4559004672, 64'd102070312, 64'd2299700480, - 64'd2391675136, - 64'd3192177152, 64'd1423954688, 64'd809671104, - 64'd3513762816, - 64'd955117760, 64'd1902938752, - 64'd631066688, - 64'd3052782592, 64'd1109274752, 64'd1558822272, - 64'd1494091520, - 64'd1556610304, 64'd2269510912, 64'd714791360, - 64'd1592675072, 64'd169091664, 64'd2305641984, - 64'd195341168, - 64'd1070712640, 64'd1423562624, 64'd1470502784, - 64'd815692352, - 64'd270500960, 64'd1848460800, 64'd283132608, - 64'd983061184, 64'd442441856, 64'd1480934400, - 64'd728544320, - 64'd742389440, 64'd821758016, 64'd646057728, - 64'd1227436800, - 64'd280649664, 64'd804295616, - 64'd233055440, - 64'd1148273920, 64'd176776304, 64'd490392160, - 64'd816879424, - 64'd657657472, 64'd459556736, 64'd67613304, - 64'd956801536, - 64'd36773232, 64'd503127744, - 64'd280112224, - 64'd705559616, 64'd451017440, 64'd347804800, - 64'd440484224, - 64'd249826912, 64'd654555200, 64'd98842528, - 64'd397910304, 64'd191381712, 64'd564903872, - 64'd128357176, - 64'd216444336, 64'd456355936, 64'd285017440, - 64'd253858800, 64'd3050629, 64'd487655872, - 64'd35300144, - 64'd254726000, 64'd169375200, 64'd328922144, - 64'd266572864, - 64'd160114736, 64'd232843824, 64'd84600728, - 64'd343313056, - 64'd28024984, 64'd194051504, - 64'd133557856, - 64'd273387424, 64'd83241808, 64'd91741472, - 64'd250064400, - 64'd117703392, 64'd136980144, - 64'd20735106, - 64'd245364816, 64'd45151444, 64'd126708256, - 64'd98853272, - 64'd149914640, 64'd152515776, 64'd71438304, - 64'd121494408, - 64'd20934352, 64'd177340880, 64'd2522624, - 64'd93310576, 64'd85350848, 64'd129883200, - 64'd51005004, - 64'd36880936, 64'd134524960, 64'd45030392, - 64'd72748896, 64'd19986240, 64'd121701616, - 64'd36592440, - 64'd62096136, 64'd55902396, 64'd66361080, - 64'd85190256, - 64'd30708068, 64'd62385892, - 64'd712312, - 64'd90387856, 64'd4752329, 64'd43981124, - 64'd51631496, - 64'd60515312, 64'd30043286, 64'd13472879, - 64'd71160592, - 64'd15059884, 64'd38102792, - 64'd14850987, - 64'd59422868, 64'd25271580, 64'd29992342, - 64'd30904236, - 64'd28217524, 64'd46593592, 64'd12575954, - 64'd31583102, 64'd6162450, 64'd45425136, - 64'd5423568, - 64'd20274662, 64'd30093992, 64'd27529158, - 64'd17130376, - 64'd4051666, 64'd37091756, 64'd3566168, - 64'd19652374, 64'd9848125, 64'd28545784, - 64'd16056442, - 64'd14220628, 64'd16770666, 64'd11336165, - 64'd25020642, - 64'd4752179, 64'd15776155, - 64'd6042734, - 64'd22494672, 64'd4252382, 64'd9111341, - 64'd17044608, - 64'd12145263, 64'd9531941, 64'd613824, - 64'd19060672, 64'd300326, 64'd9992190, - 64'd6101355, - 64'd13463918, 64'd9686351, 64'd6602173, - 64'd8942388, - 64'd4152233, 64'd13223402, 64'd1542887, - 64'd7763126, 64'd4508748, 64'd10972317, - 64'd2896221, - 64'd3957066, 64'd9430765, 64'd5146458, - 64'd5200044, 64'd428899, 64'd9656603, - 64'd1226636, - 64'd5011658, 64'd3615504, 64'd6213811, - 64'd5631469, - 64'd2991692, 64'd4693822, 64'd1260028, - 64'd6885071, - 64'd330041, 64'd3759445, - 64'd2992379, - 64'd5264326, 64'd1824922, 64'd1638819, - 64'd5117514, - 64'd2056621, 64'd2786440, - 64'd593223, - 64'd4823532, 64'd1161396, 64'd2477161, - 64'd2074662, - 64'd2793340, 64'd3182569, 64'd1313794, - 64'd2428616, - 64'd198125, 64'd3533655, - 64'd65889, - 64'd1789553, 64'd1856737, 64'd2478704, - 64'd1094159, - 64'd631857, 64'd2729918, 64'd745615, - 64'd1469285, 64'd488257, 64'd2374341, - 64'd856207, - 64'd1205504, 64'd1160352, 64'd1214091, - 64'd1758171, - 64'd552868, 64'd1238908, - 64'd125926, - 64'd1788334, 64'd152208, 64'd835064, - 64'd1101481, - 64'd1141848, 64'd633343, 64'd214239, - 64'd1433662, - 64'd220970, 64'd763440, - 64'd339770, - 64'd1150464, 64'd564573, 64'd576920, - 64'd635383, - 64'd503629, 64'd952744, 64'd218583, - 64'd623121, 64'd178576, 64'd892319, - 64'd136733, - 64'd380482, 64'd632378, 64'd512147, - 64'd356725, - 64'd52857, 64'd741974, 64'd30269, - 64'd391078, 64'd216974, 64'd547842, - 64'd348832, - 64'd270891, 64'd341680, 64'd194584, - 64'd507568, - 64'd77753, 64'd308940, - 64'd147870, - 64'd438698, 64'd98757, 64'd168294, - 64'd353873, - 64'd221901, 64'd196496, - 64'd2052, - 64'd378615, 64'd26631, 64'd197528, - 64'd131293, - 64'd255756, 64'd206340, 64'd124366, - 64'd180778, - 64'd66243, 64'd266246, 64'd21970, - 64'd150868, 64'd103193, 64'd212291, - 64'd64403, - 64'd71560, 64'd193874, 64'd91637, - 64'd106213, 64'd15757, 64'd190501, - 64'd34753, - 64'd98358, 64'd76498, 64'd116609, - 64'd118203, - 64'd55541, 64'd94217, 64'd16560, - 64'd137640, - 64'd2070, 64'd72468, - 64'd65997, - 64'd100946, 64'd39514, 64'd28739, - 64'd104297, - 64'd35151, 64'd56458, - 64'd15393, - 64'd94482, 64'd28224, 64'd48254, - 64'd43313, - 64'd51620, 64'd66025, 64'd23928, - 64'd48405, 64'd418, 64'd70157, - 64'd3596, - 64'd34171, 64'd39976, 64'd47046, - 64'd23256, - 64'd10514, 64'd55201, 64'd11795, - 64'd29554, 64'd11477, 64'd46155, - 64'd19524, - 64'd23296, 64'd23964, 64'd21972, - 64'd36118, - 64'd9799, 64'd24522, - 64'd4710, - 64'd35261, 64'd4170, 64'd15768, - 64'd23310, - 64'd21406, 64'd13271, 64'd3184, - 64'd28780, - 64'd2818, 64'd15248, - 64'd7612, - 64'd22180, 64'd12423, 64'd11048, - 64'd13002, - 64'd8839, 64'd19404, 64'd3707, - 64'd12248, 64'd4652, 64'd17468, - 64'd3283, - 64'd7087, 64'd13206, 64'd9451, - 64'd7389, - 64'd495, 64'd14791, - 64'd206, - 64'd7757, 64'd4721, 64'd10463, - 64'd7499, - 64'd5133, 64'd6935, 64'd3243, - 64'd10258, - 64'd1209, 64'd6028, - 64'd3481, - 64'd8523, 64'd2238, 64'd3079, - 64'd7310, - 64'd4008, 64'd4031, - 64'd324, - 64'd7496, 64'd938, 64'd3891, - 64'd2800, - 64'd4831, 64'd4362, 64'd2327, - 64'd3642, - 64'd989, 64'd5342, 64'd262, - 64'd2921, 64'd2314, 64'd4090, - 64'd1412, - 64'd1277, 64'd3968, 64'd1603, - 64'd2161, 64'd456, 64'd3745, - 64'd895, - 64'd1923, 64'd1607, 64'd2173, - 64'd2466, - 64'd1022, 64'd1884, 64'd160, - 64'd2742, 64'd48, 64'd1391, - 64'd1437, - 64'd1926, 64'd847, 64'd493, - 64'd2117, - 64'd583, 64'd1140, - 64'd377, - 64'd1844, 64'd661, 64'd936, - 64'd899, - 64'd945, 64'd1363, 64'd431, - 64'd962, 64'd95, 64'd1388, - 64'd117, - 64'd649, 64'd853, 64'd888, - 64'd491, - 64'd168, 64'd1112, 64'd174, - 64'd592, 64'd263, 64'd894, - 64'd437, - 64'd448, 64'd493, 64'd392, - 64'd739, - 64'd170, 64'd484, - 64'd137, - 64'd693, 64'd105, 64'd296, - 64'd490, - 64'd398, 64'd276, 64'd42, - 64'd576, - 64'd25, 64'd303, - 64'd168, - 64'd426, 64'd270, 64'd211, - 64'd265, - 64'd152, 64'd394, 64'd61, - 64'd240, 64'd114, 64'd341, - 64'd76, - 64'd131, 64'd274, 64'd173, - 64'd152, 64'd1, 64'd294, - 64'd20, - 64'd153, 64'd102, 64'd199, - 64'd160, - 64'd97, 64'd140, 64'd52, - 64'd207, - 64'd17, 64'd117, - 64'd80, - 64'd165, 64'd50, 64'd56, - 64'd150, - 64'd71, 64'd82, - 64'd12, - 64'd148, 64'd27, 64'd76, - 64'd59, - 64'd91, 64'd92, 64'd43, - 64'd73, - 64'd13, 64'd107, 64'd2, - 64'd56, 64'd51, 64'd78, - 64'd31, - 64'd22, 64'd81, 64'd27, - 64'd44, 64'd12, 64'd73, - 64'd22, - 64'd37, 64'd34, 64'd40, - 64'd51, - 64'd19, 64'd38, - 64'd0, - 64'd54, 64'd3, 64'd27, - 64'd31, - 64'd37, 64'd18, 64'd8, - 64'd43, - 64'd9, 64'd23, - 64'd9, - 64'd36, 64'd15, 64'd18, - 64'd19, - 64'd17, 64'd28, 64'd8, - 64'd19, 64'd4, 64'd27, - 64'd3, - 64'd12, 64'd18, 64'd17, - 64'd10, - 64'd2, 64'd22, 64'd2, - 64'd12, 64'd6, 64'd17, - 64'd10, - 64'd9, 64'd10, 64'd7, - 64'd15, - 64'd3, 64'd10, - 64'd4, - 64'd14, 64'd3, 64'd6, - 64'd10, - 64'd7, 64'd6, 64'd0, - 64'd11, 64'd0, 64'd6, - 64'd4, - 64'd8, 64'd6, 64'd4, - 64'd5, - 64'd3, 64'd8, 64'd1, - 64'd5, 64'd3, 64'd7, - 64'd2, - 64'd2, 64'd6, 64'd3, - 64'd3, 64'd0, 64'd6, - 64'd1, - 64'd3, 64'd2, 64'd4, - 64'd3, - 64'd2, 64'd3, 64'd1, - 64'd4, - 64'd0, 64'd2, - 64'd2, - 64'd3, 64'd1, 64'd1, - 64'd3, - 64'd1, 64'd2, - 64'd0, - 64'd3, 64'd1, 64'd1, - 64'd1, - 64'd2, 64'd2, 64'd1, - 64'd1, - 64'd0, 64'd2, - 64'd0, - 64'd1, 64'd1, 64'd1, - 64'd1, - 64'd0, 64'd2, 64'd0, - 64'd1, 64'd0, 64'd1, - 64'd1, - 64'd1, 64'd1, 64'd1, - 64'd1, - 64'd0, 64'd1, - 64'd0, - 64'd1, 64'd0, 64'd1, - 64'd1, - 64'd1, 64'd0, 64'd0, - 64'd1, - 64'd0, 64'd0, - 64'd0, - 64'd1, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd1, 64'd0, - 64'd0, 64'd0, 64'd1, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0};
	localparam logic signed[63:0] hb[0:1199] = {64'd67282986336256, 64'd15925081276416, - 64'd13053910319104, - 64'd2600907833344, 64'd46241719255040, 64'd37561451937792, - 64'd1031533821952, - 64'd5428495253504, 64'd22973836689408, 64'd42223953510400, 64'd14594550530048, - 64'd3275386781696, 64'd4008551907328, 64'd32830579015680, 64'd25656928763904, 64'd3055999516672, - 64'd6970588266496, 64'd16388061134848, 64'd27745474052096, 64'd10660821860352, - 64'd9729572077568, 64'd558183612416, 64'd21047197827072, 64'd16336497410048, - 64'd6726005817344, - 64'd9235473629184, 64'd9221060952064, 64'd18038350938112, - 64'd1572290035712, - 64'd11206951698432, - 64'd2792537194496, 64'd15519267684352, 64'd2539725258752, - 64'd6941853089792, - 64'd10944011829248, 64'd10107455799296, 64'd3868836757504, 64'd43593134080, - 64'd13410579251200, 64'd3913146171392, 64'd2363855470592, 64'd6105038061568, - 64'd10786977087488, - 64'd1098257989632, - 64'd782689632256, 64'd8878215397376, - 64'd5325878984704, - 64'd3782055559168, - 64'd3932610363392, 64'd7863339057152, 64'd265721282560, - 64'd4039707721728, - 64'd5767671840768, 64'd4165725585408, 64'd3920110813184, - 64'd2610896044032, - 64'd5743348547584, - 64'd307357745152, 64'd4809766207488, - 64'd608251281408, - 64'd4135357513728, - 64'd3761841111040, 64'd3347204800512, 64'd973607337984, - 64'd1759289540608, - 64'd5173173813248, 64'd725637267456, 64'd1587403030528, 64'd452657709056, - 64'd4498294571008, - 64'd1719660838912, 64'd1217645772800, 64'd1823868452864, - 64'd2468478976000, - 64'd3048596832256, 64'd247646093312, 64'd2125608386560, - 64'd139588567040, - 64'd2975866552320, - 64'd789078605824, 64'd1558683582464, 64'd1574487588864, - 64'd1822248665088, - 64'd1452403195904, 64'd580105928704, 64'd2206403395584, - 64'd249477169152, - 64'd1544294105088, - 64'd324482531328, 64'd1802040639488, 64'd1070292205568, - 64'd1129679159296, - 64'd825176489984, 64'd780396658688, 64'd1710814658560, - 64'd452293754880, - 64'd830565056512, - 64'd312181686272, 64'd1595238514688, 64'd197752094720, - 64'd462174879744, - 64'd1036644909056, 64'd944033038336, 64'd603327168512, 64'd44093468672, - 64'd1199774105600, 64'd123612667904, 64'd684659245056, 64'd455350353920, - 64'd867670949888, - 64'd524179013632, 64'd497407426560, 64'd629578399744, - 64'd278893756416, - 64'd803341008896, 64'd180656930816, 64'd548160176128, 64'd286385700864, - 64'd701962387456, - 64'd113976459264, 64'd294101155840, 64'd621751107584, - 64'd352735592448, - 64'd281209077760, - 64'd2937806080, 64'd654878048256, 64'd51129118720, - 64'd289786101760, - 64'd226267906048, 64'd443271741440, 64'd342598811648, - 64'd176047620096, - 64'd312955174912, 64'd122301136896, 64'd437094350848, - 64'd13857614848, - 64'd264891580416, - 64'd163707863040, 64'd344519704576, 64'd122259980288, - 64'd132998979584, - 64'd317496164352, 64'd143046770688, 64'd185387843584, 64'd13189578752, - 64'd314071711744, - 64'd66452946944, 64'd167360462848, 64'd115740844032, - 64'd192934281216, - 64'd203674533888, 64'd92692570112, 64'd147073630208, - 64'd28029116416, - 64'd234183180288, 64'd1661353472, 64'd112948879360, 64'd108060467200, - 64'd171532304384, - 64'd68537696256, 64'd42308988928, 64'd170921951232, - 64'd60893442048, - 64'd97036427264, - 64'd29120120832, 64'd154225328128, 64'd45294145536, - 64'd83297353728, - 64'd73854386176, 64'd83033202688, 64'd108645400576, - 64'd42557046784, - 64'd81010794496, - 64'd3052362496, 64'd115854442496, 64'd3562243584, - 64'd56455655424, - 64'd68188557312, 64'd77730291712, 64'd36616466432, - 64'd16636317696, - 64'd92843220992, 64'd19440162816, 64'd47458037760, 64'd20094365696, - 64'd77261340672, - 64'd32307419136, 64'd37433786368, 64'd40815644672, - 64'd36701044736, - 64'd59619008512, 64'd15378306048, 64'd41605963776, 64'd7827344896, - 64'd58019115008, - 64'd7477295104, 64'd26895316992, 64'd38786220032, - 64'd34939965440, - 64'd22283012096, 64'd5842346496, 64'd47853600768, - 64'd4111832064, - 64'd25320962048, - 64'd12203354112, 64'd36857671680, 64'd21074898944, - 64'd18181029888, - 64'd21238448128, 64'd14691079168, 64'd32507189248, - 64'd5906238976, - 64'd20055070720, - 64'd7688411648, 64'd29140660224, 64'd5716253184, - 64'd11553614848, - 64'd21846499328, 64'd15719245824, 64'd12501473280, - 64'd681912448, - 64'd24429867008, - 64'd369907456, 64'd13057359872, 64'd7902852096, - 64'd17216260096, - 64'd12487081984, 64'd8647524352, 64'd11508850688, - 64'd5232218624, - 64'd17048470528, 64'd2091785984, 64'd9951410176, 64'd5899296256, - 64'd14144353280, - 64'd3656101120, 64'd5027585536, 64'd12206102528, - 64'd6635649536, - 64'd6644591616, - 64'd626875840, 64'd12463518720, 64'd1572722304, - 64'd6416714240, - 64'd4723875840, 64'd8002545664, 64'd7240418816, - 64'd3826697984, - 64'd6098137600, 64'd1606498944, 64'd8846891008, - 64'd409438048, - 64'd4878330880, - 64'd3874911744, 64'd6752942592, 64'd2355343360, - 64'd2133099008, - 64'd6608261632, 64'd2619789312, 64'd3583894528, 64'd751143296, - 64'd6222286336, - 64'd1521067904, 64'd3177977344, 64'd2664177920, - 64'd3600797952, - 64'd4116261888, 64'd1675420032, 64'd3122017536, - 64'd254774480, - 64'd4559004672, - 64'd102070312, 64'd2299700480, 64'd2391675136, - 64'd3192177152, - 64'd1423954688, 64'd809671104, 64'd3513762816, - 64'd955117760, - 64'd1902938752, - 64'd631066688, 64'd3052782592, 64'd1109274752, - 64'd1558822272, - 64'd1494091520, 64'd1556610304, 64'd2269510912, - 64'd714791360, - 64'd1592675072, - 64'd169091664, 64'd2305641984, 64'd195341168, - 64'd1070712640, - 64'd1423562624, 64'd1470502784, 64'd815692352, - 64'd270500960, - 64'd1848460800, 64'd283132608, 64'd983061184, 64'd442441856, - 64'd1480934400, - 64'd728544320, 64'd742389440, 64'd821758016, - 64'd646057728, - 64'd1227436800, 64'd280649664, 64'd804295616, 64'd233055440, - 64'd1148273920, - 64'd176776304, 64'd490392160, 64'd816879424, - 64'd657657472, - 64'd459556736, 64'd67613304, 64'd956801536, - 64'd36773232, - 64'd503127744, - 64'd280112224, 64'd705559616, 64'd451017440, - 64'd347804800, - 64'd440484224, 64'd249826912, 64'd654555200, - 64'd98842528, - 64'd397910304, - 64'd191381712, 64'd564903872, 64'd128357176, - 64'd216444336, - 64'd456355936, 64'd285017440, 64'd253858800, 64'd3050629, - 64'd487655872, - 64'd35300144, 64'd254726000, 64'd169375200, - 64'd328922144, - 64'd266572864, 64'd160114736, 64'd232843824, - 64'd84600728, - 64'd343313056, 64'd28024984, 64'd194051504, 64'd133557856, - 64'd273387424, - 64'd83241808, 64'd91741472, 64'd250064400, - 64'd117703392, - 64'd136980144, - 64'd20735106, 64'd245364816, 64'd45151444, - 64'd126708256, - 64'd98853272, 64'd149914640, 64'd152515776, - 64'd71438304, - 64'd121494408, 64'd20934352, 64'd177340880, - 64'd2522624, - 64'd93310576, - 64'd85350848, 64'd129883200, 64'd51005004, - 64'd36880936, - 64'd134524960, 64'd45030392, 64'd72748896, 64'd19986240, - 64'd121701616, - 64'd36592440, 64'd62096136, 64'd55902396, - 64'd66361080, - 64'd85190256, 64'd30708068, 64'd62385892, 64'd712312, - 64'd90387856, - 64'd4752329, 64'd43981124, 64'd51631496, - 64'd60515312, - 64'd30043286, 64'd13472879, 64'd71160592, - 64'd15059884, - 64'd38102792, - 64'd14850987, 64'd59422868, 64'd25271580, - 64'd29992342, - 64'd30904236, 64'd28217524, 64'd46593592, - 64'd12575954, - 64'd31583102, - 64'd6162450, 64'd45425136, 64'd5423568, - 64'd20274662, - 64'd30093992, 64'd27529158, 64'd17130376, - 64'd4051666, - 64'd37091756, 64'd3566168, 64'd19652374, 64'd9848125, - 64'd28545784, - 64'd16056442, 64'd14220628, 64'd16770666, - 64'd11336165, - 64'd25020642, 64'd4752179, 64'd15776155, 64'd6042734, - 64'd22494672, - 64'd4252382, 64'd9111341, 64'd17044608, - 64'd12145263, - 64'd9531941, 64'd613824, 64'd19060672, 64'd300326, - 64'd9992190, - 64'd6101355, 64'd13463918, 64'd9686351, - 64'd6602173, - 64'd8942388, 64'd4152233, 64'd13223402, - 64'd1542887, - 64'd7763126, - 64'd4508748, 64'd10972317, 64'd2896221, - 64'd3957066, - 64'd9430765, 64'd5146458, 64'd5200044, 64'd428899, - 64'd9656603, - 64'd1226636, 64'd5011658, 64'd3615504, - 64'd6213811, - 64'd5631469, 64'd2991692, 64'd4693822, - 64'd1260028, - 64'd6885071, 64'd330041, 64'd3759445, 64'd2992379, - 64'd5264326, - 64'd1824922, 64'd1638819, 64'd5117514, - 64'd2056621, - 64'd2786440, - 64'd593223, 64'd4823532, 64'd1161396, - 64'd2477161, - 64'd2074662, 64'd2793340, 64'd3182569, - 64'd1313794, - 64'd2428616, 64'd198125, 64'd3533655, 64'd65889, - 64'd1789553, - 64'd1856737, 64'd2478704, 64'd1094159, - 64'd631857, - 64'd2729918, 64'd745615, 64'd1469285, 64'd488257, - 64'd2374341, - 64'd856207, 64'd1205504, 64'd1160352, - 64'd1214091, - 64'd1758171, 64'd552868, 64'd1238908, 64'd125926, - 64'd1788334, - 64'd152208, 64'd835064, 64'd1101481, - 64'd1141848, - 64'd633343, 64'd214239, 64'd1433662, - 64'd220970, - 64'd763440, - 64'd339770, 64'd1150464, 64'd564573, - 64'd576920, - 64'd635383, 64'd503629, 64'd952744, - 64'd218583, - 64'd623121, - 64'd178576, 64'd892319, 64'd136733, - 64'd380482, - 64'd632378, 64'd512147, 64'd356725, - 64'd52857, - 64'd741974, 64'd30269, 64'd391078, 64'd216974, - 64'd547842, - 64'd348832, 64'd270891, 64'd341680, - 64'd194584, - 64'd507568, 64'd77753, 64'd308940, 64'd147870, - 64'd438698, - 64'd98757, 64'd168294, 64'd353873, - 64'd221901, - 64'd196496, - 64'd2052, 64'd378615, 64'd26631, - 64'd197528, - 64'd131293, 64'd255756, 64'd206340, - 64'd124366, - 64'd180778, 64'd66243, 64'd266246, - 64'd21970, - 64'd150868, - 64'd103193, 64'd212291, 64'd64403, - 64'd71560, - 64'd193874, 64'd91637, 64'd106213, 64'd15757, - 64'd190501, - 64'd34753, 64'd98358, 64'd76498, - 64'd116609, - 64'd118203, 64'd55541, 64'd94217, - 64'd16560, - 64'd137640, 64'd2070, 64'd72468, 64'd65997, - 64'd100946, - 64'd39514, 64'd28739, 64'd104297, - 64'd35151, - 64'd56458, - 64'd15393, 64'd94482, 64'd28224, - 64'd48254, - 64'd43313, 64'd51620, 64'd66025, - 64'd23928, - 64'd48405, - 64'd418, 64'd70157, 64'd3596, - 64'd34171, - 64'd39976, 64'd47046, 64'd23256, - 64'd10514, - 64'd55201, 64'd11795, 64'd29554, 64'd11477, - 64'd46155, - 64'd19524, 64'd23296, 64'd23964, - 64'd21972, - 64'd36118, 64'd9799, 64'd24522, 64'd4710, - 64'd35261, - 64'd4170, 64'd15768, 64'd23310, - 64'd21406, - 64'd13271, 64'd3184, 64'd28780, - 64'd2818, - 64'd15248, - 64'd7612, 64'd22180, 64'd12423, - 64'd11048, - 64'd13002, 64'd8839, 64'd19404, - 64'd3707, - 64'd12248, - 64'd4652, 64'd17468, 64'd3283, - 64'd7087, - 64'd13206, 64'd9451, 64'd7389, - 64'd495, - 64'd14791, - 64'd206, 64'd7757, 64'd4721, - 64'd10463, - 64'd7499, 64'd5133, 64'd6935, - 64'd3243, - 64'd10258, 64'd1209, 64'd6028, 64'd3481, - 64'd8523, - 64'd2238, 64'd3079, 64'd7310, - 64'd4008, - 64'd4031, - 64'd324, 64'd7496, 64'd938, - 64'd3891, - 64'd2800, 64'd4831, 64'd4362, - 64'd2327, - 64'd3642, 64'd989, 64'd5342, - 64'd262, - 64'd2921, - 64'd2314, 64'd4090, 64'd1412, - 64'd1277, - 64'd3968, 64'd1603, 64'd2161, 64'd456, - 64'd3745, - 64'd895, 64'd1923, 64'd1607, - 64'd2173, - 64'd2466, 64'd1022, 64'd1884, - 64'd160, - 64'd2742, - 64'd48, 64'd1391, 64'd1437, - 64'd1926, - 64'd847, 64'd493, 64'd2117, - 64'd583, - 64'd1140, - 64'd377, 64'd1844, 64'd661, - 64'd936, - 64'd899, 64'd945, 64'd1363, - 64'd431, - 64'd962, - 64'd95, 64'd1388, 64'd117, - 64'd649, - 64'd853, 64'd888, 64'd491, - 64'd168, - 64'd1112, 64'd174, 64'd592, 64'd263, - 64'd894, - 64'd437, 64'd448, 64'd493, - 64'd392, - 64'd739, 64'd170, 64'd484, 64'd137, - 64'd693, - 64'd105, 64'd296, 64'd490, - 64'd398, - 64'd276, 64'd42, 64'd576, - 64'd25, - 64'd303, - 64'd168, 64'd426, 64'd270, - 64'd211, - 64'd265, 64'd152, 64'd394, - 64'd61, - 64'd240, - 64'd114, 64'd341, 64'd76, - 64'd131, - 64'd274, 64'd173, 64'd152, 64'd1, - 64'd294, - 64'd20, 64'd153, 64'd102, - 64'd199, - 64'd160, 64'd97, 64'd140, - 64'd52, - 64'd207, 64'd17, 64'd117, 64'd80, - 64'd165, - 64'd50, 64'd56, 64'd150, - 64'd71, - 64'd82, - 64'd12, 64'd148, 64'd27, - 64'd76, - 64'd59, 64'd91, 64'd92, - 64'd43, - 64'd73, 64'd13, 64'd107, - 64'd2, - 64'd56, - 64'd51, 64'd78, 64'd31, - 64'd22, - 64'd81, 64'd27, 64'd44, 64'd12, - 64'd73, - 64'd22, 64'd37, 64'd34, - 64'd40, - 64'd51, 64'd19, 64'd38, 64'd0, - 64'd54, - 64'd3, 64'd27, 64'd31, - 64'd37, - 64'd18, 64'd8, 64'd43, - 64'd9, - 64'd23, - 64'd9, 64'd36, 64'd15, - 64'd18, - 64'd19, 64'd17, 64'd28, - 64'd8, - 64'd19, - 64'd4, 64'd27, 64'd3, - 64'd12, - 64'd18, 64'd17, 64'd10, - 64'd2, - 64'd22, 64'd2, 64'd12, 64'd6, - 64'd17, - 64'd10, 64'd9, 64'd10, - 64'd7, - 64'd15, 64'd3, 64'd10, 64'd4, - 64'd14, - 64'd3, 64'd6, 64'd10, - 64'd7, - 64'd6, 64'd0, 64'd11, 64'd0, - 64'd6, - 64'd4, 64'd8, 64'd6, - 64'd4, - 64'd5, 64'd3, 64'd8, - 64'd1, - 64'd5, - 64'd3, 64'd7, 64'd2, - 64'd2, - 64'd6, 64'd3, 64'd3, 64'd0, - 64'd6, - 64'd1, 64'd3, 64'd2, - 64'd4, - 64'd3, 64'd2, 64'd3, - 64'd1, - 64'd4, 64'd0, 64'd2, 64'd2, - 64'd3, - 64'd1, 64'd1, 64'd3, - 64'd1, - 64'd2, - 64'd0, 64'd3, 64'd1, - 64'd1, - 64'd1, 64'd2, 64'd2, - 64'd1, - 64'd1, 64'd0, 64'd2, 64'd0, - 64'd1, - 64'd1, 64'd1, 64'd1, - 64'd0, - 64'd2, 64'd0, 64'd1, 64'd0, - 64'd1, - 64'd1, 64'd1, 64'd1, - 64'd1, - 64'd1, 64'd0, 64'd1, 64'd0, - 64'd1, - 64'd0, 64'd1, 64'd1, - 64'd1, - 64'd0, 64'd0, 64'd1, - 64'd0, - 64'd0, - 64'd0, 64'd1, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd1, - 64'd0, - 64'd0, - 64'd0, 64'd1, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0, 64'd0, 64'd0, 64'd0, - 64'd0, - 64'd0};
endpackage
`endif
