
module LUT #(
    parameter       size = 1,
    parameter real  re[size-1:0],
                    im[size-1:0]
) (
    input logic[size-1:0] sel,
    output complex result
);
    // Generate LUT values
    complex mem[2**size-1:0];
    genvar i;
    generate
        for(i = 0; i < size**2; i++) begin
            mem[i].r = rtof(calcLUT(size, re, j));
            mem[i].i = rtof(calcLUT(size, im, j));
        end
    endgenerate

    always_comb begin : select
        result = mem[sel];
    end
endmodule

function real calcLUT(int size, real fact[size-1:0], logic[size-1:0] in);
    real temp = 0.0;
    logic[size:0] j;
    for(j = 0; j < size; j++) begin
        if(in[j] == 1) begin
            temp += fact[j];
        end else begin
            temp -= fact[j];
        end
    end
    calcLUT = temp;
endfunction