`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam N = 3;
	localparam M = 3;
	localparam real Lfr[0:2] = {0.92746544, 0.9558213, 0.9558213};
	localparam real Lfi[0:2] = {0.0, 0.10899793, -0.10899793};
	localparam real Lbr[0:2] = {0.92746544, 0.9558213, 0.9558213};
	localparam real Lbi[0:2] = {0.0, 0.10899793, -0.10899793};
	localparam real Wfr[0:2] = {-0.0024392875, 0.001540601, 0.001540601};
	localparam real Wfi[0:2] = {-0.0, -0.0028816545, 0.0028816545};
	localparam real Wbr[0:2] = {0.0024392875, -0.001540601, -0.001540601};
	localparam real Wbi[0:2] = {0.0, 0.0028816545, -0.0028816545};
	localparam real Ffr[0:2][0:74] = '{
		'{-8.178999, 1.2289, -0.33600852, -7.5857387, 1.1397622, -0.3116363, -7.0355105, 1.05709, -0.2890319, -6.5251927, 0.9804145, -0.2680671, -6.051891, 0.90930057, -0.24862297, -5.61292, 0.84334487, -0.23058921, -5.205789, 0.7821732, -0.21386352, -4.8281894, 0.7254386, -0.19835103, -4.4779787, 0.67281926, -0.18396373, -4.1531706, 0.6240166, -0.17062, -3.8519223, 0.5787538, -0.15824415, -3.5725248, 0.53677416, -0.14676598, -3.3133934, 0.4978395, -0.13612038, -3.0730577, 0.46172893, -0.12624694, -2.8501549, 0.42823762, -0.11708968, -2.6434202, 0.3971756, -0.10859663, -2.451681, 0.36836666, -0.10071962, -2.2738492, 0.34164733, -0.09341397, -2.1089165, 0.3168661, -0.08663823, -1.9559473, 0.29388237, -0.08035396, -1.8140736, 0.27256572, -0.07452552, -1.6824905, 0.2527953, -0.06911985, -1.5604517, 0.2344589, -0.06410627, -1.4472651, 0.21745253, -0.059456352, -1.3422884, 0.2016797, -0.05514371},
		'{4.244545, -0.69897884, -0.06948673, 3.879046, -0.7595571, -0.045866925, 3.4871297, -0.8051144, -0.023372946, 3.076186, -0.8361399, -0.002232031, 2.6533172, -0.8532875, 0.017364228, 2.2252612, -0.8573543, 0.035259888, 1.7983255, -0.8492587, 0.051334146, 1.3783324, -0.8300193, 0.06550039, 0.97057384, -0.8007326, 0.077704884, 0.5797782, -0.76255256, 0.087924995, 0.21008697, -0.71667004, 0.096167244, -0.13495895, -0.66429365, 0.102465026, -0.45242348, -0.60663193, 0.106876135, -0.73997086, -0.54487634, 0.109480165, -0.99585325, -0.48018622, 0.11037576, -1.218891, -0.41367504, 0.109677866, -1.4084468, -0.34639853, 0.10751488, -1.5643939, -0.27934432, 0.104025915, -1.6870798, -0.21342336, 0.099358045, -1.7772863, -0.14946301, 0.0936637, -1.8361862, -0.08820191, 0.08709814, -1.8652979, -0.030286266, 0.07981711, -1.8664386, 0.02373214, 0.07197464, -1.8416772, 0.07339655, 0.06372107, -1.7932866, 0.11834447, 0.055201177},
		'{4.244545, -0.69897884, -0.06948673, 3.879046, -0.7595571, -0.045866925, 3.4871297, -0.8051144, -0.023372946, 3.076186, -0.8361399, -0.002232031, 2.6533172, -0.8532875, 0.017364228, 2.2252612, -0.8573543, 0.035259888, 1.7983255, -0.8492587, 0.051334146, 1.3783324, -0.8300193, 0.06550039, 0.97057384, -0.8007326, 0.077704884, 0.5797782, -0.76255256, 0.087924995, 0.21008697, -0.71667004, 0.096167244, -0.13495895, -0.66429365, 0.102465026, -0.45242348, -0.60663193, 0.106876135, -0.73997086, -0.54487634, 0.109480165, -0.99585325, -0.48018622, 0.11037576, -1.218891, -0.41367504, 0.109677866, -1.4084468, -0.34639853, 0.10751488, -1.5643939, -0.27934432, 0.104025915, -1.6870798, -0.21342336, 0.099358045, -1.7772863, -0.14946301, 0.0936637, -1.8361862, -0.08820191, 0.08709814, -1.8652979, -0.030286266, 0.07981711, -1.8664386, 0.02373214, 0.07197464, -1.8416772, 0.07339655, 0.06372107, -1.7932866, 0.11834447, 0.055201177}};
	localparam real Ffi[0:2][0:74] = '{
		'{0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0},
		'{1.6328791, 0.8390828, -0.18853539, 2.0233872, 0.7258259, -0.18778005, 2.3568046, 0.6109697, -0.18448357, 2.6327739, 0.49622205, -0.17888093, 2.8517592, 0.38316208, -0.1712215, 3.0149782, 0.2732279, -0.16176449, 3.1243293, 0.1677072, -0.15077469, 3.1823142, 0.06773068, -0.13851833, 3.1919591, -0.025731964, -0.12525937, 3.156733, -0.11187336, -0.1112559, 3.0804672, -0.19004759, -0.096757114, 2.9672751, -0.2597671, -0.08200048, 2.8214746, -0.32069755, -0.067209326, 2.6475122, -0.37265116, -0.05259083, 2.4498932, -0.4155783, -0.03833432, 2.2331142, -0.4495579, -0.02461003, 2.0016015, -0.47478673, -0.011568131, 1.7596555, -0.491568, 0.00066183356, 1.5114005, -0.5002991, 0.011971204, 1.2607405, -0.50145924, 0.022272153, 1.0113221, -0.4955966, 0.031497348, 0.76650274, -0.4833156, 0.03959935, 0.529326, -0.46526447, 0.0465498, 0.30250314, -0.44212294, 0.05233838, 0.088399924, -0.41459045, 0.056971602},
		'{-1.6328791, -0.8390828, 0.18853539, -2.0233872, -0.7258259, 0.18778005, -2.3568046, -0.6109697, 0.18448357, -2.6327739, -0.49622205, 0.17888093, -2.8517592, -0.38316208, 0.1712215, -3.0149782, -0.2732279, 0.16176449, -3.1243293, -0.1677072, 0.15077469, -3.1823142, -0.06773068, 0.13851833, -3.1919591, 0.025731964, 0.12525937, -3.156733, 0.11187336, 0.1112559, -3.0804672, 0.19004759, 0.096757114, -2.9672751, 0.2597671, 0.08200048, -2.8214746, 0.32069755, 0.067209326, -2.6475122, 0.37265116, 0.05259083, -2.4498932, 0.4155783, 0.03833432, -2.2331142, 0.4495579, 0.02461003, -2.0016015, 0.47478673, 0.011568131, -1.7596555, 0.491568, -0.00066183356, -1.5114005, 0.5002991, -0.011971204, -1.2607405, 0.50145924, -0.022272153, -1.0113221, 0.4955966, -0.031497348, -0.76650274, 0.4833156, -0.03959935, -0.529326, 0.46526447, -0.0465498, -0.30250314, 0.44212294, -0.05233838, -0.088399924, 0.41459045, -0.056971602}};
	localparam real Fbr[0:2][0:74] = '{
		'{8.178999, 1.2289, 0.33600852, 7.5857387, 1.1397622, 0.3116363, 7.0355105, 1.05709, 0.2890319, 6.5251927, 0.9804145, 0.2680671, 6.051891, 0.90930057, 0.24862297, 5.61292, 0.84334487, 0.23058921, 5.205789, 0.7821732, 0.21386352, 4.8281894, 0.7254386, 0.19835103, 4.4779787, 0.67281926, 0.18396373, 4.1531706, 0.6240166, 0.17062, 3.8519223, 0.5787538, 0.15824415, 3.5725248, 0.53677416, 0.14676598, 3.3133934, 0.4978395, 0.13612038, 3.0730577, 0.46172893, 0.12624694, 2.8501549, 0.42823762, 0.11708968, 2.6434202, 0.3971756, 0.10859663, 2.451681, 0.36836666, 0.10071962, 2.2738492, 0.34164733, 0.09341397, 2.1089165, 0.3168661, 0.08663823, 1.9559473, 0.29388237, 0.08035396, 1.8140736, 0.27256572, 0.07452552, 1.6824905, 0.2527953, 0.06911985, 1.5604517, 0.2344589, 0.06410627, 1.4472651, 0.21745253, 0.059456352, 1.3422884, 0.2016797, 0.05514371},
		'{-4.244545, -0.69897884, 0.06948673, -3.879046, -0.7595571, 0.045866925, -3.4871297, -0.8051144, 0.023372946, -3.076186, -0.8361399, 0.002232031, -2.6533172, -0.8532875, -0.017364228, -2.2252612, -0.8573543, -0.035259888, -1.7983255, -0.8492587, -0.051334146, -1.3783324, -0.8300193, -0.06550039, -0.97057384, -0.8007326, -0.077704884, -0.5797782, -0.76255256, -0.087924995, -0.21008697, -0.71667004, -0.096167244, 0.13495895, -0.66429365, -0.102465026, 0.45242348, -0.60663193, -0.106876135, 0.73997086, -0.54487634, -0.109480165, 0.99585325, -0.48018622, -0.11037576, 1.218891, -0.41367504, -0.109677866, 1.4084468, -0.34639853, -0.10751488, 1.5643939, -0.27934432, -0.104025915, 1.6870798, -0.21342336, -0.099358045, 1.7772863, -0.14946301, -0.0936637, 1.8361862, -0.08820191, -0.08709814, 1.8652979, -0.030286266, -0.07981711, 1.8664386, 0.02373214, -0.07197464, 1.8416772, 0.07339655, -0.06372107, 1.7932866, 0.11834447, -0.055201177},
		'{-4.244545, -0.69897884, 0.06948673, -3.879046, -0.7595571, 0.045866925, -3.4871297, -0.8051144, 0.023372946, -3.076186, -0.8361399, 0.002232031, -2.6533172, -0.8532875, -0.017364228, -2.2252612, -0.8573543, -0.035259888, -1.7983255, -0.8492587, -0.051334146, -1.3783324, -0.8300193, -0.06550039, -0.97057384, -0.8007326, -0.077704884, -0.5797782, -0.76255256, -0.087924995, -0.21008697, -0.71667004, -0.096167244, 0.13495895, -0.66429365, -0.102465026, 0.45242348, -0.60663193, -0.106876135, 0.73997086, -0.54487634, -0.109480165, 0.99585325, -0.48018622, -0.11037576, 1.218891, -0.41367504, -0.109677866, 1.4084468, -0.34639853, -0.10751488, 1.5643939, -0.27934432, -0.104025915, 1.6870798, -0.21342336, -0.099358045, 1.7772863, -0.14946301, -0.0936637, 1.8361862, -0.08820191, -0.08709814, 1.8652979, -0.030286266, -0.07981711, 1.8664386, 0.02373214, -0.07197464, 1.8416772, 0.07339655, -0.06372107, 1.7932866, 0.11834447, -0.055201177}};
	localparam real Fbi[0:2][0:74] = '{
		'{0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0},
		'{-1.6328791, 0.8390828, 0.18853539, -2.0233872, 0.7258259, 0.18778005, -2.3568046, 0.6109697, 0.18448357, -2.6327739, 0.49622205, 0.17888093, -2.8517592, 0.38316208, 0.1712215, -3.0149782, 0.2732279, 0.16176449, -3.1243293, 0.1677072, 0.15077469, -3.1823142, 0.06773068, 0.13851833, -3.1919591, -0.025731964, 0.12525937, -3.156733, -0.11187336, 0.1112559, -3.0804672, -0.19004759, 0.096757114, -2.9672751, -0.2597671, 0.08200048, -2.8214746, -0.32069755, 0.067209326, -2.6475122, -0.37265116, 0.05259083, -2.4498932, -0.4155783, 0.03833432, -2.2331142, -0.4495579, 0.02461003, -2.0016015, -0.47478673, 0.011568131, -1.7596555, -0.491568, -0.00066183356, -1.5114005, -0.5002991, -0.011971204, -1.2607405, -0.50145924, -0.022272153, -1.0113221, -0.4955966, -0.031497348, -0.76650274, -0.4833156, -0.03959935, -0.529326, -0.46526447, -0.0465498, -0.30250314, -0.44212294, -0.05233838, -0.088399924, -0.41459045, -0.056971602},
		'{1.6328791, -0.8390828, -0.18853539, 2.0233872, -0.7258259, -0.18778005, 2.3568046, -0.6109697, -0.18448357, 2.6327739, -0.49622205, -0.17888093, 2.8517592, -0.38316208, -0.1712215, 3.0149782, -0.2732279, -0.16176449, 3.1243293, -0.1677072, -0.15077469, 3.1823142, -0.06773068, -0.13851833, 3.1919591, 0.025731964, -0.12525937, 3.156733, 0.11187336, -0.1112559, 3.0804672, 0.19004759, -0.096757114, 2.9672751, 0.2597671, -0.08200048, 2.8214746, 0.32069755, -0.067209326, 2.6475122, 0.37265116, -0.05259083, 2.4498932, 0.4155783, -0.03833432, 2.2331142, 0.4495579, -0.02461003, 2.0016015, 0.47478673, -0.011568131, 1.7596555, 0.491568, 0.00066183356, 1.5114005, 0.5002991, 0.011971204, 1.2607405, 0.50145924, 0.022272153, 1.0113221, 0.4955966, 0.031497348, 0.76650274, 0.4833156, 0.03959935, 0.529326, 0.46526447, 0.0465498, 0.30250314, 0.44212294, 0.05233838, 0.088399924, 0.41459045, 0.056971602}};
	localparam real hf[0:899] = {0.042440016, -0.00031544187, -0.00048106903, 0.042117327, -0.00093739753, -0.00046338927, 0.041489176, -0.0015380593, -0.00043022074, 0.04056866, -0.0021079478, -0.00038393072, 0.03937328, -0.002638915, -0.00032683677, 0.037924256, -0.0031241453, -0.0002611825, 0.036245894, -0.0035581344, -0.00018911558, 0.034364924, -0.0039366577, -0.00011266883, 0.032309856, -0.0042567197, -3.374357e-05, 0.030110419, -0.004516495, 4.5903784e-05, 0.02779695, -0.004715255, 0.00012467254, 0.025399903, -0.0048532872, 0.00020112577, 0.02294934, -0.0049318084, 0.00027399557, 0.020474503, -0.0049528675, 0.0003421859, 0.018003413, -0.0049192514, 0.00040477287, 0.015562539, -0.004834383, 0.00046100284, 0.013176492, -0.004702219, 0.00051028846, 0.010867797, -0.0045271507, 0.00055220275, 0.008656688, -0.004313906, 0.0005864715, 0.0065609766, -0.004067454, 0.0006129645, 0.004595948, -0.0037929101, 0.0006316851, 0.0027743103, -0.0034954555, 0.0006427591, 0.0011061853, -0.003180252, 0.0006464229, -0.000400865, -0.0028523707, 0.00064301083, -0.0017417748, -0.0025167244, 0.00063294225, -0.00291388, -0.0021780082, 0.00061670865, -0.003916796, -0.0018406484, 0.0005948606, -0.0047522713, -0.0015087576, 0.0005679949, -0.005424022, -0.0011860991, 0.0005367424, -0.0059375498, -0.00087605877, 0.0005017558, -0.0062999455, -0.0005816237, 0.00046369867, -0.006519689, -0.00030536868, 0.00042323463, -0.006606439, -4.9449438e-05, 0.00038101783, -0.006570825, 0.00018439768, 0.00033768412, -0.006424236, 0.00039485015, 0.00029384304, -0.0061786207, 0.00058098824, 0.00025007108, -0.0058462853, 0.00074227905, 0.00020690575, -0.005439709, 0.0008785566, 0.00016484059, -0.0049713636, 0.0009899975, 0.00012432142, -0.0044535515, 0.0010770947, 8.574336e-05, -0.0038982537, 0.0011406278, 4.9448885e-05, -0.0033169948, 0.0011816317, 1.5726711e-05, -0.002720723, 0.0012013646, -1.5188404e-05, -0.002119708, 0.0012012743, -4.3115127e-05, -0.0015234547, 0.0011829654, -6.792429e-05, -0.000940632, 0.0011481654, -8.953696e-05, -0.0003790215, 0.0010986931, -0.00010792201, 0.00015452123, 0.0010364266, -0.00012309312, 0.0006540881, 0.00096327387, -0.00013510541, 0.0011147262, 0.00088114425, -0.00014405174, 0.001532432, 0.000791923, -0.00015005877, 0.0019041329, 0.00069744705, -0.00015328276, 0.0022276572, 0.00059948367, -0.00015390536, 0.002501695, 0.0004997117, -0.0001521293, 0.0027257493, 0.0003997054, -0.00014817412, 0.00290008, 0.00030092036, -0.00014227194, 0.0030256421, 0.00020468306, -0.00013466344, 0.003104019, 0.00011218207, -0.00012559396, 0.0031373505, 2.446228e-05, -0.00011530983, 0.0031282625, -5.7578578e-05, -0.00010405493, 0.0030797906, -0.00013319119, -9.206762e-05, 0.0029953076, -0.00020177376, -7.957784e-05, 0.00287845, -0.00026286909, -6.6804685e-05, 0.0027330467, -0.00031615997, -5.3954176e-05, 0.0025630502, -0.000361463, -4.1217467e-05, 0.002372473, -0.00039872093, -2.8769331e-05, 0.0021653248, -0.00042799397, -1.676701e-05, 0.0019455578, -0.00044945, -5.34939e-06, 0.0017170149, -0.00046335414, 5.3635254e-06, 0.0014833839, -0.00047005774, 1.5270833e-05, 0.0012481575, -0.0004699869, 2.4290674e-05, 0.0010145985, -0.00046363103, 3.2359912e-05, 0.0007857118, -0.00045153112, 3.9433606e-05, 0.0005642207, -0.00043426844, 4.548422e-05, 0.0003525504, -0.0004124534, 5.0500712e-05, 0.00015281576, -0.00038671485, 5.448743e-05, -3.3185224e-05, -0.00035768986, 5.7462883e-05, -0.00020397302, -0.0003260144, 5.9458405e-05, -0.00035838372, -0.00029231436, 6.051677e-05, -0.00049556204, -0.0002571978, 6.069071e-05, -0.0006149504, -0.00022124762, 6.004144e-05, -0.0007162748, -0.0001850155, 5.8637175e-05, -0.00079952774, -0.00014901638, 5.6551635e-05, -0.000864949, -0.000113724236, 5.3862615e-05, -0.0009130037, -7.956831e-05, 5.0650593e-05, -0.0009443595, -4.6930665e-05, 4.6997407e-05, -0.0009598628, -1.6144268e-05, 4.2985008e-05, -0.0009605132, 1.2507932e-05, 3.8694317e-05, -0.0009474392, 3.879324e-05, 3.4204175e-05, -0.0009218728, 6.2528714e-05, 2.9590388e-05, -0.0008851248, 8.358e-05, 2.4924917e-05, -0.00083856116, 0.000101859616, 2.0275147e-05, -0.00078357995, 0.00011732464, 1.57033e-05, -0.00072159007, 0.00012997408, 1.1265945e-05, -0.0006539906, 0.0001398457, 7.0136443e-06, -0.0005821527, 0.00014701266, 2.9906848e-06, -0.0005074026, 0.00015157992, -7.6506353e-07, -0.00043100672, 0.00015368036, -4.2222e-06, -0.0003541589, 0.00015347093, -7.355749e-06, -0.00027796908, 0.00015112867, -1.0147028e-05, -0.00020345443, 0.00014684678, -1.2583442e-05, -0.0001315323, 0.00014083077, -1.4658207e-05, -6.301494e-05, 0.00013329467, -1.6370013e-05, 1.3937813e-06, 0.0001244575, -1.7722636e-05, 6.11e-05, 0.000114539835, -1.872451e-05, 0.00011561982, 0.00010376065, -1.9388262e-05, 0.00016457777, 9.2334434e-05, -1.9730236e-05, 0.00020770384, 8.0468555e-05, -1.9769981e-05, 0.00024482937, 6.8360925e-05, -1.9529745e-05, 0.00027588176, 5.6197976e-05, -1.903398e-05, 0.00030087825, 4.4152956e-05, -1.8308821e-05, 0.000319919, 3.238449e-05, -1.7381617e-05, 0.0003331795, 2.1035505e-05, -1.6280459e-05, 0.00034090245, 1.0232421e-05, -1.503373e-05, 0.0003433894, 8.463261e-08, -1.3669702e-05, 0.00034099218, -9.3157305e-06, -1.2216148e-05, 0.00033410423, -1.7893784e-05, -1.0699999e-05, 0.00032315208, -2.559164e-05, -9.14703e-06, 0.00030858692, -3.236794e-05, -7.5816006e-06, 0.00029087655, -3.8197188e-05, -6.026412e-06, 0.00027049755, -4.3068914e-05, -4.502326e-06, 0.0002479282, -4.6986715e-05, -3.0282108e-06, 0.00022364152, -4.9967133e-05, -1.6208293e-06, 0.00019809927, -5.203847e-05, -2.9476516e-07, 0.00017174632, -5.3239528e-05, 9.3761577e-07, 0.0001450057, -5.361826e-05, 2.0661714e-06, 0.00011827447, -5.323045e-05, 3.0829572e-06, 9.192005e-05, -5.213835e-05, 3.982172e-06, 6.6277404e-05, -5.0409326e-05, 4.760078e-06, 4.1646792e-05, -4.8114554e-05, 5.4148977e-06, 1.8292207e-05, -4.5327743e-05, 5.9466943e-06, -3.5596015e-06, -4.2123927e-05, 6.3572306e-06, -2.3719474e-05, -3.8578342e-05, 6.6498196e-06, -4.2035677e-05, -3.4765337e-05, 6.8291615e-06, -5.8393205e-05, -3.075745e-05, 6.901176e-06, -7.271265e-05, -2.6624502e-05, 6.87283e-06, -8.494866e-05, -2.2432863e-05, 6.7519604e-06, -9.5088006e-05, -1.8244771e-05, 6.5471036e-06, -0.0001031474, -1.4117787e-05, 6.267323e-06, -0.00010917102, -1.0104344e-05, 5.922046e-06, -0.00011322788, -6.2514036e-06, 5.5209043e-06, -0.00011540899, -2.6002156e-06, 5.0735866e-06, -0.0001158245, 8.138305e-07, 4.5897004e-06, -0.00011460072, 3.961256e-06, 4.0786445e-06, -0.000111877205, 6.818462e-06, 3.5494943e-06, -0.00010780381, 9.367619e-06, 3.0109002e-06, -0.000102537866, 1.159648e-05, 2.4710005e-06, -9.624145e-05, 1.3498141e-05, 1.9373454e-06, -8.907878e-05, 1.507073e-05, 1.4168379e-06, -8.1213795e-05, 1.6317066e-05, 9.156852e-07, -7.280792e-05, 1.7244267e-05, 4.3936518e-07, -6.401799e-05, 1.786333e-05, -7.3950397e-09, -5.4994474e-05, 1.8188694e-05, -4.2062882e-07, -4.5879817e-05, 1.8237779e-05, -7.9712817e-07, -3.68071e-05, 1.803053e-05, -1.1344315e-06, -2.789889e-05, 1.7588944e-05, -1.4308023e-06, -1.9266332e-05, 1.6936623e-05, -1.6851991e-06, -1.10084575e-05, 1.6098318e-05, -1.897238e-06, -3.2117266e-06, 1.509951e-05, -2.0671494e-06, 4.050235e-06, 1.3965999e-05, -2.195728e-06, 1.0716697e-05, 1.2723521e-05, -2.2842817e-06, 1.6739701e-05, 1.1397404e-05, -2.3345735e-06, 2.2083774e-05, 1.001224e-05, -2.3487637e-06, 2.6725484e-05, 8.591607e-06, -2.3293512e-06, 3.065287e-05, 7.157814e-06, -2.2791126e-06, 3.386475e-05, 5.7316875e-06, -2.2010443e-06, 3.6369933e-05, 4.3323957e-06, -2.0983032e-06, 3.8186354e-05, 2.9773068e-06, -1.9741528e-06, 3.9340142e-05, 1.6818814e-06, -1.831909e-06, 3.986466e-05, 4.5960175e-07, -1.6748904e-06, 3.9799474e-05, -6.780666e-07, -1.5063728e-06, 3.918938e-05, -1.7216839e-06, -1.3295463e-06, 3.8083374e-05, -2.6638156e-06, -1.1474785e-06, 3.6533656e-05, -3.4989853e-06, -9.630805e-07, 3.459469e-05, -4.223605e-06, -7.790785e-07, 3.232226e-05, -4.835884e-06, -5.9798987e-07, 2.9772604e-05, -5.335719e-06, -4.2210414e-07, 2.7001617e-05, -5.72457e-06, -2.5346793e-07, 2.406409e-05, -6.005325e-06, -9.387508e-08, 2.1013031e-05, -6.182151e-06, 5.513954e-08, 1.7899076e-05, -6.260343e-06, 1.9230183e-07, 1.4769958e-05, -6.246166e-06, 3.1659664e-07, 1.1670065e-05, -6.146696e-06, 4.2726265e-07, 8.640072e-06, -5.9696617e-06, 5.2378374e-07, 5.7166603e-06, -5.7232896e-06, 6.0587803e-07, 2.932304e-06, -5.4161515e-06, 6.7348435e-07, 3.1513457e-07, -5.057021e-06, 7.2674646e-07, -2.1111234e-06, -4.654739e-06, 7.659959e-07, -4.327153e-06, -4.2180823e-06, 7.917333e-07, -6.3179846e-06, -3.755651e-06, 8.0460916e-07, -8.072877e-06, -3.2757603e-06, 8.0540326e-07, -9.585152e-06, -2.786347e-06, 7.950044e-07, -1.0851985e-05, -2.2948893e-06, 7.743902e-07, -1.18741555e-05, -1.8083352e-06, 7.446065e-07, -1.2655769e-05, -1.3330483e-06, 7.0674827e-07, -1.320395e-05, -8.747616e-07, 6.619406e-07, -1.3528523e-05, -4.3854604e-07, 6.1132073e-07, -1.3641669e-05, -2.8789307e-08, 5.560217e-07, -1.3557589e-05, 3.5081365e-07, 4.971568e-07, -1.3292151e-05, 6.9726036e-07, 4.358058e-07, -1.286255e-05, 1.0082307e-06, 3.7300225e-07, -1.2286966e-05, 1.2820678e-06, 3.0972288e-07, -1.1584249e-05, 1.5177525e-06, 2.4687824e-07, -1.0773596e-05, 1.7148684e-06, 1.8530497e-07, -9.874271e-06, 1.8735643e-06, 1.2575984e-07, -8.905327e-06, 1.994509e-06, 6.891516e-08, -7.885358e-06, 2.0788432e-06, 1.53558e-08, -6.8322797e-06, 2.1281298e-06, -3.4422392e-08, -5.763129e-06, 2.1442995e-06, -8.001282e-08, -4.693897e-06, 2.129597e-06, -1.2109707e-07, -3.6393824e-06, 2.086527e-06, -1.5744284e-07, -2.6130774e-06, 2.0177997e-06, -1.889006e-07, -1.6270786e-06, 1.9262784e-06, -2.1539964e-07, -6.9202343e-07, 1.814928e-06, -2.3694304e-07, 1.8294848e-07, 1.6867671e-06, -2.5360225e-07, 9.902099e-07, 1.5448212e-06, -2.655109e-07, 1.7236384e-06, 1.3920817e-06, -2.7285836e-07, 2.37859e-06, 1.2314658e-06, -2.7588302e-07, 2.9518515e-06, 1.0657826e-06, -2.748653e-07, 3.44158e-06, 8.977016e-07, -2.7012055e-07, 3.8472253e-06, 7.2972676e-07, -2.6199226e-07, 4.169441e-06, 5.641739e-07, -2.5084503e-07, 4.409987e-06, 4.0315257e-07, -2.3705815e-07, 4.571621e-06, 2.4855262e-07, -2.2101905e-07, 4.657987e-06, 1.0203409e-07, -2.0311748e-07, 4.673499e-06, -3.4978427e-08, -1.8373993e-07, 4.6232212e-06, -1.6129805e-07, -1.6326445e-07, 4.5127517e-06, -2.7597423e-07, -1.4205611e-07, 4.3481036e-06, -3.7828832e-07, -1.2046296e-07, 4.1355916e-06, -4.677463e-07, -9.881236e-08, 3.8817207e-06, -5.440687e-07, -7.74081e-08, 3.5930846e-06, -6.071787e-07, -5.6527934e-08, 3.2762662e-06, -6.571879e-07, -3.642164e-08, 2.9377472e-06, -6.9438073e-07, -1.730968e-08, 2.5838274e-06, -7.1919794e-07, 6.1765787e-10, 2.2205493e-06, -7.322183e-07, 1.7200666e-08, 1.8536348e-06, -7.34141e-07, 3.231013e-08, 1.4884298e-06, -7.2576626e-07, 4.584685e-08, 1.1298582e-06, -7.079774e-07, 5.7740777e-08, 7.823851e-07, -6.8172193e-07, 6.7949806e-08, 4.4998947e-07, -6.47994e-07, 7.645827e-08, 1.3614515e-07, -6.0781696e-07, 8.3275204e-08, -1.5618951e-07, -5.6222717e-07, 8.8432365e-08, -4.245741e-07, -5.1225857e-07, 9.198211e-08, -6.670814e-07, -4.589286e-07, 9.39951e-08, -8.8228563e-07, -4.0322547e-07, 9.4558025e-08, -1.0692451e-06, -3.460965e-07, 9.377115e-08, -1.2274787e-06, -2.884381e-07, 9.1745946e-08, -1.3569389e-06, -2.3108728e-07, 8.860271e-08, -1.4579794e-06, -1.7481439e-07, 8.446823e-08, -1.5313204e-06, -1.2031745e-07, 7.947356e-08, -1.5780124e-06, -6.82179e-08, 7.375189e-08, -1.5993953e-06, -1.9057726e-08, 6.7436545e-08, -1.5970597e-06, 2.6702159e-08, 6.065911e-08, -1.5728058e-06, 6.868221e-08, 5.3547765e-08, -1.5286025e-06, 1.06583464e-07, 4.6225765e-08, -1.4665482e-06, 1.4018563e-07, 3.8810075e-08, -1.3888315e-06, 1.6934433e-07, 3.141026e-08, -1.2976948e-06, 1.9398739e-07, 2.412748e-08, -1.195399e-06, 2.1411049e-07, 1.7053756e-08, -1.0841908e-06, 2.2977213e-07, 1.02713456e-08, -9.662726e-07, 2.4108817e-07, 3.8523544e-09, -8.4377575e-07, 2.4822594e-07, -2.141515e-09, -7.1873586e-07, 2.5139815e-07, -7.659039e-09, -5.930722e-07, 2.508564e-07, -1.2659397e-08, -4.6856934e-07, 2.4688504e-07, -1.7111969e-08, -3.4686312e-07, 2.3979456e-07, -2.099599e-08, -2.2942862e-07, 2.2991549e-07, -2.4300109e-08, -1.1757191e-07, 2.1759232e-07, -2.702184e-08, -1.2424563e-08, 2.0317766e-07, -2.916694e-08, 8.505896e-08, 1.8702679e-07, -3.0748716e-08, 1.7410136e-07, 1.6949248e-07, -3.1787263e-08, 2.541e-07, 1.5092039e-07, -3.2308705e-08, 3.246223e-07, 1.3164477e-07, -3.234437e-08, 3.8539898e-07, 1.1198465e-07, -3.1929968e-08, 4.363156e-07, 9.224066e-08, -3.1104772e-08, 4.7740264e-07, 7.2692146e-08, -2.9910808e-08, 5.0882437e-07, 5.3594956e-08, -2.8392082e-08, 5.3086643e-07, 3.5179603e-08, -2.6593801e-08, 5.439229e-07, 1.7650011e-08, -2.4561674e-08, 5.484829e-07, 1.1826409e-09, -2.2341236e-08, 5.451164e-07, -1.4073883e-08, -1.9977241e-08, 5.3446075e-07, -2.7998766e-08, -1.7513083e-08, 5.1720656e-07, -4.049863e-08, -1.4990313e-08, 4.9408425e-07, -5.1506778e-08, -1.2448197e-08, 4.6585092e-07, -6.09821e-08, -9.923339e-09, 4.3327802e-07, -6.8907774e-08, -7.449378e-09, 3.9713953e-07, -7.528965e-08, -5.0567426e-09, 3.58201e-07, -8.01545e-08, -2.7724674e-09, 3.1720973e-07, -8.3548095e-08, -6.2007416e-10, 2.748857e-07, -8.553313e-08, 1.3804927e-09, 2.3191366e-07, -8.618713e-08, 3.2128753e-09, 1.889363e-07, -8.560023e-08, 4.8642614e-09, 1.4654847e-07, -8.387303e-08, 6.325297e-09, 1.05292585e-07, -8.111441e-08, 7.589958e-09, 6.5654916e-08, -7.743938e-08, 8.655387e-09, 2.8063155e-08, -7.2967076e-08, 9.521692e-09, -7.1151978e-09, -6.781878e-08, 1.0191732e-08, -3.9573408e-08, -6.211608e-08, 1.0670863e-08, -6.906522e-08, -5.5979168e-08, 1.0966687e-08};
	localparam real hb[0:899] = {0.042440016, 0.00031544187, -0.00048106903, 0.042117327, 0.00093739753, -0.00046338927, 0.041489176, 0.0015380593, -0.00043022074, 0.04056866, 0.0021079478, -0.00038393072, 0.03937328, 0.002638915, -0.00032683677, 0.037924256, 0.0031241453, -0.0002611825, 0.036245894, 0.0035581344, -0.00018911558, 0.034364924, 0.0039366577, -0.00011266883, 0.032309856, 0.0042567197, -3.374357e-05, 0.030110419, 0.004516495, 4.5903784e-05, 0.02779695, 0.004715255, 0.00012467254, 0.025399903, 0.0048532872, 0.00020112577, 0.02294934, 0.0049318084, 0.00027399557, 0.020474503, 0.0049528675, 0.0003421859, 0.018003413, 0.0049192514, 0.00040477287, 0.015562539, 0.004834383, 0.00046100284, 0.013176492, 0.004702219, 0.00051028846, 0.010867797, 0.0045271507, 0.00055220275, 0.008656688, 0.004313906, 0.0005864715, 0.0065609766, 0.004067454, 0.0006129645, 0.004595948, 0.0037929101, 0.0006316851, 0.0027743103, 0.0034954555, 0.0006427591, 0.0011061853, 0.003180252, 0.0006464229, -0.000400865, 0.0028523707, 0.00064301083, -0.0017417748, 0.0025167244, 0.00063294225, -0.00291388, 0.0021780082, 0.00061670865, -0.003916796, 0.0018406484, 0.0005948606, -0.0047522713, 0.0015087576, 0.0005679949, -0.005424022, 0.0011860991, 0.0005367424, -0.0059375498, 0.00087605877, 0.0005017558, -0.0062999455, 0.0005816237, 0.00046369867, -0.006519689, 0.00030536868, 0.00042323463, -0.006606439, 4.9449438e-05, 0.00038101783, -0.006570825, -0.00018439768, 0.00033768412, -0.006424236, -0.00039485015, 0.00029384304, -0.0061786207, -0.00058098824, 0.00025007108, -0.0058462853, -0.00074227905, 0.00020690575, -0.005439709, -0.0008785566, 0.00016484059, -0.0049713636, -0.0009899975, 0.00012432142, -0.0044535515, -0.0010770947, 8.574336e-05, -0.0038982537, -0.0011406278, 4.9448885e-05, -0.0033169948, -0.0011816317, 1.5726711e-05, -0.002720723, -0.0012013646, -1.5188404e-05, -0.002119708, -0.0012012743, -4.3115127e-05, -0.0015234547, -0.0011829654, -6.792429e-05, -0.000940632, -0.0011481654, -8.953696e-05, -0.0003790215, -0.0010986931, -0.00010792201, 0.00015452123, -0.0010364266, -0.00012309312, 0.0006540881, -0.00096327387, -0.00013510541, 0.0011147262, -0.00088114425, -0.00014405174, 0.001532432, -0.000791923, -0.00015005877, 0.0019041329, -0.00069744705, -0.00015328276, 0.0022276572, -0.00059948367, -0.00015390536, 0.002501695, -0.0004997117, -0.0001521293, 0.0027257493, -0.0003997054, -0.00014817412, 0.00290008, -0.00030092036, -0.00014227194, 0.0030256421, -0.00020468306, -0.00013466344, 0.003104019, -0.00011218207, -0.00012559396, 0.0031373505, -2.446228e-05, -0.00011530983, 0.0031282625, 5.7578578e-05, -0.00010405493, 0.0030797906, 0.00013319119, -9.206762e-05, 0.0029953076, 0.00020177376, -7.957784e-05, 0.00287845, 0.00026286909, -6.6804685e-05, 0.0027330467, 0.00031615997, -5.3954176e-05, 0.0025630502, 0.000361463, -4.1217467e-05, 0.002372473, 0.00039872093, -2.8769331e-05, 0.0021653248, 0.00042799397, -1.676701e-05, 0.0019455578, 0.00044945, -5.34939e-06, 0.0017170149, 0.00046335414, 5.3635254e-06, 0.0014833839, 0.00047005774, 1.5270833e-05, 0.0012481575, 0.0004699869, 2.4290674e-05, 0.0010145985, 0.00046363103, 3.2359912e-05, 0.0007857118, 0.00045153112, 3.9433606e-05, 0.0005642207, 0.00043426844, 4.548422e-05, 0.0003525504, 0.0004124534, 5.0500712e-05, 0.00015281576, 0.00038671485, 5.448743e-05, -3.3185224e-05, 0.00035768986, 5.7462883e-05, -0.00020397302, 0.0003260144, 5.9458405e-05, -0.00035838372, 0.00029231436, 6.051677e-05, -0.00049556204, 0.0002571978, 6.069071e-05, -0.0006149504, 0.00022124762, 6.004144e-05, -0.0007162748, 0.0001850155, 5.8637175e-05, -0.00079952774, 0.00014901638, 5.6551635e-05, -0.000864949, 0.000113724236, 5.3862615e-05, -0.0009130037, 7.956831e-05, 5.0650593e-05, -0.0009443595, 4.6930665e-05, 4.6997407e-05, -0.0009598628, 1.6144268e-05, 4.2985008e-05, -0.0009605132, -1.2507932e-05, 3.8694317e-05, -0.0009474392, -3.879324e-05, 3.4204175e-05, -0.0009218728, -6.2528714e-05, 2.9590388e-05, -0.0008851248, -8.358e-05, 2.4924917e-05, -0.00083856116, -0.000101859616, 2.0275147e-05, -0.00078357995, -0.00011732464, 1.57033e-05, -0.00072159007, -0.00012997408, 1.1265945e-05, -0.0006539906, -0.0001398457, 7.0136443e-06, -0.0005821527, -0.00014701266, 2.9906848e-06, -0.0005074026, -0.00015157992, -7.6506353e-07, -0.00043100672, -0.00015368036, -4.2222e-06, -0.0003541589, -0.00015347093, -7.355749e-06, -0.00027796908, -0.00015112867, -1.0147028e-05, -0.00020345443, -0.00014684678, -1.2583442e-05, -0.0001315323, -0.00014083077, -1.4658207e-05, -6.301494e-05, -0.00013329467, -1.6370013e-05, 1.3937813e-06, -0.0001244575, -1.7722636e-05, 6.11e-05, -0.000114539835, -1.872451e-05, 0.00011561982, -0.00010376065, -1.9388262e-05, 0.00016457777, -9.2334434e-05, -1.9730236e-05, 0.00020770384, -8.0468555e-05, -1.9769981e-05, 0.00024482937, -6.8360925e-05, -1.9529745e-05, 0.00027588176, -5.6197976e-05, -1.903398e-05, 0.00030087825, -4.4152956e-05, -1.8308821e-05, 0.000319919, -3.238449e-05, -1.7381617e-05, 0.0003331795, -2.1035505e-05, -1.6280459e-05, 0.00034090245, -1.0232421e-05, -1.503373e-05, 0.0003433894, -8.463261e-08, -1.3669702e-05, 0.00034099218, 9.3157305e-06, -1.2216148e-05, 0.00033410423, 1.7893784e-05, -1.0699999e-05, 0.00032315208, 2.559164e-05, -9.14703e-06, 0.00030858692, 3.236794e-05, -7.5816006e-06, 0.00029087655, 3.8197188e-05, -6.026412e-06, 0.00027049755, 4.3068914e-05, -4.502326e-06, 0.0002479282, 4.6986715e-05, -3.0282108e-06, 0.00022364152, 4.9967133e-05, -1.6208293e-06, 0.00019809927, 5.203847e-05, -2.9476516e-07, 0.00017174632, 5.3239528e-05, 9.3761577e-07, 0.0001450057, 5.361826e-05, 2.0661714e-06, 0.00011827447, 5.323045e-05, 3.0829572e-06, 9.192005e-05, 5.213835e-05, 3.982172e-06, 6.6277404e-05, 5.0409326e-05, 4.760078e-06, 4.1646792e-05, 4.8114554e-05, 5.4148977e-06, 1.8292207e-05, 4.5327743e-05, 5.9466943e-06, -3.5596015e-06, 4.2123927e-05, 6.3572306e-06, -2.3719474e-05, 3.8578342e-05, 6.6498196e-06, -4.2035677e-05, 3.4765337e-05, 6.8291615e-06, -5.8393205e-05, 3.075745e-05, 6.901176e-06, -7.271265e-05, 2.6624502e-05, 6.87283e-06, -8.494866e-05, 2.2432863e-05, 6.7519604e-06, -9.5088006e-05, 1.8244771e-05, 6.5471036e-06, -0.0001031474, 1.4117787e-05, 6.267323e-06, -0.00010917102, 1.0104344e-05, 5.922046e-06, -0.00011322788, 6.2514036e-06, 5.5209043e-06, -0.00011540899, 2.6002156e-06, 5.0735866e-06, -0.0001158245, -8.138305e-07, 4.5897004e-06, -0.00011460072, -3.961256e-06, 4.0786445e-06, -0.000111877205, -6.818462e-06, 3.5494943e-06, -0.00010780381, -9.367619e-06, 3.0109002e-06, -0.000102537866, -1.159648e-05, 2.4710005e-06, -9.624145e-05, -1.3498141e-05, 1.9373454e-06, -8.907878e-05, -1.507073e-05, 1.4168379e-06, -8.1213795e-05, -1.6317066e-05, 9.156852e-07, -7.280792e-05, -1.7244267e-05, 4.3936518e-07, -6.401799e-05, -1.786333e-05, -7.3950397e-09, -5.4994474e-05, -1.8188694e-05, -4.2062882e-07, -4.5879817e-05, -1.8237779e-05, -7.9712817e-07, -3.68071e-05, -1.803053e-05, -1.1344315e-06, -2.789889e-05, -1.7588944e-05, -1.4308023e-06, -1.9266332e-05, -1.6936623e-05, -1.6851991e-06, -1.10084575e-05, -1.6098318e-05, -1.897238e-06, -3.2117266e-06, -1.509951e-05, -2.0671494e-06, 4.050235e-06, -1.3965999e-05, -2.195728e-06, 1.0716697e-05, -1.2723521e-05, -2.2842817e-06, 1.6739701e-05, -1.1397404e-05, -2.3345735e-06, 2.2083774e-05, -1.001224e-05, -2.3487637e-06, 2.6725484e-05, -8.591607e-06, -2.3293512e-06, 3.065287e-05, -7.157814e-06, -2.2791126e-06, 3.386475e-05, -5.7316875e-06, -2.2010443e-06, 3.6369933e-05, -4.3323957e-06, -2.0983032e-06, 3.8186354e-05, -2.9773068e-06, -1.9741528e-06, 3.9340142e-05, -1.6818814e-06, -1.831909e-06, 3.986466e-05, -4.5960175e-07, -1.6748904e-06, 3.9799474e-05, 6.780666e-07, -1.5063728e-06, 3.918938e-05, 1.7216839e-06, -1.3295463e-06, 3.8083374e-05, 2.6638156e-06, -1.1474785e-06, 3.6533656e-05, 3.4989853e-06, -9.630805e-07, 3.459469e-05, 4.223605e-06, -7.790785e-07, 3.232226e-05, 4.835884e-06, -5.9798987e-07, 2.9772604e-05, 5.335719e-06, -4.2210414e-07, 2.7001617e-05, 5.72457e-06, -2.5346793e-07, 2.406409e-05, 6.005325e-06, -9.387508e-08, 2.1013031e-05, 6.182151e-06, 5.513954e-08, 1.7899076e-05, 6.260343e-06, 1.9230183e-07, 1.4769958e-05, 6.246166e-06, 3.1659664e-07, 1.1670065e-05, 6.146696e-06, 4.2726265e-07, 8.640072e-06, 5.9696617e-06, 5.2378374e-07, 5.7166603e-06, 5.7232896e-06, 6.0587803e-07, 2.932304e-06, 5.4161515e-06, 6.7348435e-07, 3.1513457e-07, 5.057021e-06, 7.2674646e-07, -2.1111234e-06, 4.654739e-06, 7.659959e-07, -4.327153e-06, 4.2180823e-06, 7.917333e-07, -6.3179846e-06, 3.755651e-06, 8.0460916e-07, -8.072877e-06, 3.2757603e-06, 8.0540326e-07, -9.585152e-06, 2.786347e-06, 7.950044e-07, -1.0851985e-05, 2.2948893e-06, 7.743902e-07, -1.18741555e-05, 1.8083352e-06, 7.446065e-07, -1.2655769e-05, 1.3330483e-06, 7.0674827e-07, -1.320395e-05, 8.747616e-07, 6.619406e-07, -1.3528523e-05, 4.3854604e-07, 6.1132073e-07, -1.3641669e-05, 2.8789307e-08, 5.560217e-07, -1.3557589e-05, -3.5081365e-07, 4.971568e-07, -1.3292151e-05, -6.9726036e-07, 4.358058e-07, -1.286255e-05, -1.0082307e-06, 3.7300225e-07, -1.2286966e-05, -1.2820678e-06, 3.0972288e-07, -1.1584249e-05, -1.5177525e-06, 2.4687824e-07, -1.0773596e-05, -1.7148684e-06, 1.8530497e-07, -9.874271e-06, -1.8735643e-06, 1.2575984e-07, -8.905327e-06, -1.994509e-06, 6.891516e-08, -7.885358e-06, -2.0788432e-06, 1.53558e-08, -6.8322797e-06, -2.1281298e-06, -3.4422392e-08, -5.763129e-06, -2.1442995e-06, -8.001282e-08, -4.693897e-06, -2.129597e-06, -1.2109707e-07, -3.6393824e-06, -2.086527e-06, -1.5744284e-07, -2.6130774e-06, -2.0177997e-06, -1.889006e-07, -1.6270786e-06, -1.9262784e-06, -2.1539964e-07, -6.9202343e-07, -1.814928e-06, -2.3694304e-07, 1.8294848e-07, -1.6867671e-06, -2.5360225e-07, 9.902099e-07, -1.5448212e-06, -2.655109e-07, 1.7236384e-06, -1.3920817e-06, -2.7285836e-07, 2.37859e-06, -1.2314658e-06, -2.7588302e-07, 2.9518515e-06, -1.0657826e-06, -2.748653e-07, 3.44158e-06, -8.977016e-07, -2.7012055e-07, 3.8472253e-06, -7.2972676e-07, -2.6199226e-07, 4.169441e-06, -5.641739e-07, -2.5084503e-07, 4.409987e-06, -4.0315257e-07, -2.3705815e-07, 4.571621e-06, -2.4855262e-07, -2.2101905e-07, 4.657987e-06, -1.0203409e-07, -2.0311748e-07, 4.673499e-06, 3.4978427e-08, -1.8373993e-07, 4.6232212e-06, 1.6129805e-07, -1.6326445e-07, 4.5127517e-06, 2.7597423e-07, -1.4205611e-07, 4.3481036e-06, 3.7828832e-07, -1.2046296e-07, 4.1355916e-06, 4.677463e-07, -9.881236e-08, 3.8817207e-06, 5.440687e-07, -7.74081e-08, 3.5930846e-06, 6.071787e-07, -5.6527934e-08, 3.2762662e-06, 6.571879e-07, -3.642164e-08, 2.9377472e-06, 6.9438073e-07, -1.730968e-08, 2.5838274e-06, 7.1919794e-07, 6.1765787e-10, 2.2205493e-06, 7.322183e-07, 1.7200666e-08, 1.8536348e-06, 7.34141e-07, 3.231013e-08, 1.4884298e-06, 7.2576626e-07, 4.584685e-08, 1.1298582e-06, 7.079774e-07, 5.7740777e-08, 7.823851e-07, 6.8172193e-07, 6.7949806e-08, 4.4998947e-07, 6.47994e-07, 7.645827e-08, 1.3614515e-07, 6.0781696e-07, 8.3275204e-08, -1.5618951e-07, 5.6222717e-07, 8.8432365e-08, -4.245741e-07, 5.1225857e-07, 9.198211e-08, -6.670814e-07, 4.589286e-07, 9.39951e-08, -8.8228563e-07, 4.0322547e-07, 9.4558025e-08, -1.0692451e-06, 3.460965e-07, 9.377115e-08, -1.2274787e-06, 2.884381e-07, 9.1745946e-08, -1.3569389e-06, 2.3108728e-07, 8.860271e-08, -1.4579794e-06, 1.7481439e-07, 8.446823e-08, -1.5313204e-06, 1.2031745e-07, 7.947356e-08, -1.5780124e-06, 6.82179e-08, 7.375189e-08, -1.5993953e-06, 1.9057726e-08, 6.7436545e-08, -1.5970597e-06, -2.6702159e-08, 6.065911e-08, -1.5728058e-06, -6.868221e-08, 5.3547765e-08, -1.5286025e-06, -1.06583464e-07, 4.6225765e-08, -1.4665482e-06, -1.4018563e-07, 3.8810075e-08, -1.3888315e-06, -1.6934433e-07, 3.141026e-08, -1.2976948e-06, -1.9398739e-07, 2.412748e-08, -1.195399e-06, -2.1411049e-07, 1.7053756e-08, -1.0841908e-06, -2.2977213e-07, 1.02713456e-08, -9.662726e-07, -2.4108817e-07, 3.8523544e-09, -8.4377575e-07, -2.4822594e-07, -2.141515e-09, -7.1873586e-07, -2.5139815e-07, -7.659039e-09, -5.930722e-07, -2.508564e-07, -1.2659397e-08, -4.6856934e-07, -2.4688504e-07, -1.7111969e-08, -3.4686312e-07, -2.3979456e-07, -2.099599e-08, -2.2942862e-07, -2.2991549e-07, -2.4300109e-08, -1.1757191e-07, -2.1759232e-07, -2.702184e-08, -1.2424563e-08, -2.0317766e-07, -2.916694e-08, 8.505896e-08, -1.8702679e-07, -3.0748716e-08, 1.7410136e-07, -1.6949248e-07, -3.1787263e-08, 2.541e-07, -1.5092039e-07, -3.2308705e-08, 3.246223e-07, -1.3164477e-07, -3.234437e-08, 3.8539898e-07, -1.1198465e-07, -3.1929968e-08, 4.363156e-07, -9.224066e-08, -3.1104772e-08, 4.7740264e-07, -7.2692146e-08, -2.9910808e-08, 5.0882437e-07, -5.3594956e-08, -2.8392082e-08, 5.3086643e-07, -3.5179603e-08, -2.6593801e-08, 5.439229e-07, -1.7650011e-08, -2.4561674e-08, 5.484829e-07, -1.1826409e-09, -2.2341236e-08, 5.451164e-07, 1.4073883e-08, -1.9977241e-08, 5.3446075e-07, 2.7998766e-08, -1.7513083e-08, 5.1720656e-07, 4.049863e-08, -1.4990313e-08, 4.9408425e-07, 5.1506778e-08, -1.2448197e-08, 4.6585092e-07, 6.09821e-08, -9.923339e-09, 4.3327802e-07, 6.8907774e-08, -7.449378e-09, 3.9713953e-07, 7.528965e-08, -5.0567426e-09, 3.58201e-07, 8.01545e-08, -2.7724674e-09, 3.1720973e-07, 8.3548095e-08, -6.2007416e-10, 2.748857e-07, 8.553313e-08, 1.3804927e-09, 2.3191366e-07, 8.618713e-08, 3.2128753e-09, 1.889363e-07, 8.560023e-08, 4.8642614e-09, 1.4654847e-07, 8.387303e-08, 6.325297e-09, 1.05292585e-07, 8.111441e-08, 7.589958e-09, 6.5654916e-08, 7.743938e-08, 8.655387e-09, 2.8063155e-08, 7.2967076e-08, 9.521692e-09, -7.1151978e-09, 6.781878e-08, 1.0191732e-08, -3.9573408e-08, 6.211608e-08, 1.0670863e-08, -6.906522e-08, 5.5979168e-08, 1.0966687e-08};
endpackage
`endif
