`ifndef data/Coefficients_SV_
`define data/Coefficients_SV_
package data/Coefficients;
	localparam N = 4;
	localparam real Lfr[0:3] = {0.9858421395544803, 0.9858421395544803, 0.9781171130721753, 0.9781171130721753};
	localparam real Lfi[0:3] = {0.10665246939093465, -0.10665246939093465, 0.04106261390834118, -0.04106261390834118};
	localparam real Lbr[0:3] = {0.9858421395544803, 0.9858421395544803, 0.9781171130721753, 0.9781171130721753};
	localparam real Lbi[0:3] = {0.10665246939093465, -0.10665246939093465, 0.04106261390834118, -0.04106261390834118};
	localparam real Wfr[0:3] = {8.595154768326466e-05, 8.595154768326466e-05, -2.802177544383421e-05, -2.802177544383421e-05};
	localparam real Wfi[0:3] = {0.00010408412209034592, -0.00010408412209034592, -0.00011768972452177725, 0.00011768972452177725};
	localparam real Wbr[0:3] = {-8.595154768326466e-05, -8.595154768326466e-05, 2.802177544383421e-05, 2.802177544383421e-05};
	localparam real Wbi[0:3] = {-0.00010408412209034592, 0.00010408412209034592, 0.00011768972452177725, -0.00011768972452177725};
	localparam real Ffr[0:3][0:79] = '{
		'{9.517403442589092, 5.803958733344014, -0.4775028600506327, -0.051475557707039, 12.334175399393775, 5.453185696094708, -0.5490632879926326, -0.04322707994592666, 14.96102263415146, 5.045163100567296, -0.6130702424751429, -0.03461632419982426, 17.37071831975333, 4.585572275315287, -0.6689092796911043, -0.025749026363305512, 19.53900499187631, 4.080596352735773, -0.7160707871752784, -0.01673212178091013, 21.444825625147537, 3.5368402976503113, -0.7541541277356487, -0.007672487370335698, 23.070513795269598, 2.9612473918572286, -0.7828704526032709, 0.0013242945205483789, 24.401941410865636, 2.3610132006917723, -0.8020441735158046, 0.010155136578104976, 25.428623015324696, 1.7434980596004206, -0.8116130991452264, 0.018720598010421204, 26.143776178374335, 1.1161391184899858, -0.8116272566501304, 0.02692597454909598, 26.544338013417295, 0.486362969358328, -0.802246434005084, 0.03468231537764404, 26.630938363918823, -0.1385001412055984, -0.7837364929699213, 0.04190735643865942, 26.407830694600133, -0.7512995481769507, -0.7564645159572013, 0.048526360716390216, 25.882782195429897, -1.345143932141644, -0.7208928624949469, 0.05447285732557144, 25.066925053280514, -1.913476746075026, -0.677572222336209, 0.05968927254545548, 23.974571262882375, -2.4501465043811197, -0.6271337624237217, 0.06412744730359313, 22.622993731046726, -2.949471206591621, -0.5702804737794054, 0.06774903702028089, 21.03217677218664, -3.406296248196691, -0.5077778318738266, 0.0705257911547416, 19.224539395604726, -3.8160452573072905, -0.4404438900763632, 0.07243971123109369, 17.224635043031086, -4.174763387130108, -0.36913893034683815, 0.0734830875492399},
		'{9.51740344258746, 5.803958733344131, -0.47750286005066395, -0.05147555770703265, 12.334175399392215, 5.45318569609482, -0.5490632879926624, -0.043227079945920587, 14.961022634149993, 5.045163100567405, -0.613070242475171, -0.03461632419981855, 17.37071831975197, 4.585572275315388, -0.6689092796911302, -0.0257490263633002, 19.53900499187507, 4.080596352735866, -0.716070787175302, -0.016732121780905287, 21.444825625146432, 3.5368402976503965, -0.7541541277356698, -0.0076724873703313615, 23.07051379526864, 2.961247391857304, -0.7828704526032892, 0.0013242945205521675, 24.401941410864822, 2.361013200691838, -0.8020441735158201, 0.010155136578108175, 25.428623015324046, 1.743498059600476, -0.8116130991452388, 0.018720598010423785, 26.143776178373848, 1.1161391184900298, -0.8116272566501396, 0.026925974549097925, 26.544338013416983, 0.4863629693583609, -0.8022464340050901, 0.03468231537764534, 26.63093836391867, -0.1385001412055773, -0.7837364929699241, 0.041907356438660066, 26.407830694600147, -0.7512995481769416, -0.7564645159572009, 0.04852636071639022, 25.882782195430078, -1.3451439321416463, -0.7208928624949434, 0.054472857325570806, 25.06692505328085, -1.9134767460750393, -0.6775722223362024, 0.05968927254545422, 23.974571262882865, -2.450146504381144, -0.6271337624237122, 0.0641274473035913, 22.62299373104736, -2.949471206591656, -0.5702804737793931, 0.06774903702027849, 21.032176772187412, -3.406296248196736, -0.507777831873812, 0.07052579115473867, 19.224539395605618, -3.8160452573073442, -0.44044389007634605, 0.07243971123109028, 17.224635043032087, -4.17476338713017, -0.3691389303468188, 0.07348308754923608},
		'{-9.313313592773765, -5.688953814066472, 0.40599510904134345, -0.19382811981932202, -12.087015729293103, -5.405857783345071, 0.3589502986526131, -0.18671439091601966, -14.719161330735629, -5.1228350901578645, 0.31308546179083796, -0.17949236217734052, -17.209940666047885, -4.8404954274546945, 0.2684508079689891, -0.17218217464535937, -19.559842146665797, -4.559421645725951, 0.22509179460033948, -0.16480332234289366, -21.769638866145826, -4.280169607798952, 0.18304922627424028, -0.1573746369854663, -23.840375083421378, -4.003268108103177, 0.14235935997530536, -0.14991427476315658, -25.77335268129348, -3.7292188538971804, 0.10305401577095727, -0.14243970513484921, -27.570117630503294, -3.4584965059201647, 0.0651606925002054, -0.13496770157542248, -29.23244648845956, -3.191548775908135, 0.0287026880051382, -0.1275143342146665, -30.762332960409537, -2.9287965783978374, -0.006300776544155451, -0.12009496430516839, -32.16197454955081, -2.6706342342314704, -0.039834428670685595, -0.11272424045505701, -33.43375932128638, -2.417429723170744, -0.07188681338676661, -0.10541609656034238, -34.58025280553011, -2.169524983030432, -0.10245015918354083, -0.09818375137062299, -35.60418505967578, -1.927236252748512, -0.13152024162071368, -0.09103970962115071, -36.508437913554964, -1.6908544568223671, -0.15909624491166258, -0.0839957646636417, -37.2960324164273, -1.4606456285578837, -0.18518062188698006, -0.07706300252778789, -37.9701165047758, -1.2368513696004657, -0.2097789527070889, -0.07025180734515825, -38.53395290842061, -1.0196893432437162, -0.23289980268185642, -0.06357186806706984, -38.990907311220546, -0.8093537990426116, -0.2545545795421773, -0.05703218640805522},
		'{-9.313313592769488, -5.688953814066671, 0.40599510904141745, -0.1938281198193366, -12.08701572928894, -5.405857783345265, 0.35895029865268496, -0.18671439091603384, -14.71916133073158, -5.122835090158053, 0.31308546179090785, -0.1794923621773543, -17.209940666043956, -4.8404954274548775, 0.2684508079690569, -0.17218217464537272, -19.559842146661993, -4.559421645726127, 0.22509179460040502, -0.1648033223429066, -21.769638866142145, -4.280169607799123, 0.18304922627430356, -0.15737463698547874, -23.84037508341783, -4.0032681081033425, 0.14235935997536636, -0.14991427476316863, -25.773352681290067, -3.729218853897339, 0.10305401577101594, -0.14243970513486076, -27.570117630500015, -3.4584965059203165, 0.06516069250026163, -0.13496770157543359, -29.232446488456414, -3.191548775908281, 0.0287026880051921, -0.12751433421467714, -30.76233296040653, -2.9287965783979777, -0.0063007765441039365, -0.12009496430517856, -32.161974549547935, -2.6706342342316036, -0.039834428670636524, -0.1127242404550667, -33.43375932128365, -2.41742972317087, -0.07188681338671998, -0.10541609656035161, -34.580252805527515, -2.169524983030552, -0.10245015918349654, -0.09818375137063172, -35.60418505967332, -1.9272362527486258, -0.13152024162067183, -0.09103970962115898, -36.50843791355265, -1.6908544568224744, -0.1590962449116232, -0.0839957646636495, -37.29603241642513, -1.4606456285579843, -0.1851806218869431, -0.0770630025277952, -37.97011650477375, -1.23685136960056, -0.2097789527070543, -0.0702518073451651, -38.5339529084187, -1.0196893432438041, -0.23289980268182417, -0.06357186806707624, -38.99090731121877, -0.8093537990426936, -0.25455457954214733, -0.05703218640806115}};
	localparam real Ffi[0:3][0:79] = '{
		'{-27.674164915298654, 2.5184733274811264, 0.7343556810658382, -0.07050651561734925, -26.267303371139647, 3.101823664729105, 0.6730319166502996, -0.07499828955147023, -24.57994429148466, 3.639504198693084, 0.6049442691826638, -0.07854674905514027, -22.636314861901248, 4.12605570931263, 0.5309940973721856, -0.08112661160071676, -20.463203071189568, 4.556702195122724, 0.4521355305666279, -0.08272422960131473, -18.089604766013927, 4.927394718959295, 0.3693635411114507, -0.0833375536092401, -15.546351057642116, 5.234846103754052, 0.2837017436183584, -0.08297596187978651, -12.865720722547834, 5.476556229982367, 0.1961900669407216, -0.08165996051034236, -10.081042334625243, 5.650827799274608, 0.10787244368610588, -0.07942075979239319, -7.226290906310707, 5.756772541325502, 0.01978465946861291, -0.07629973375248889, -4.335683799492918, 5.794307952239594, -0.06705750012583211, -0.0723477710935723, -1.4432805958451844, 5.764144760575793, -0.15166967264393882, -0.06762452686766418, 1.4174085081242387, 5.667765421397218, -0.2331097869118613, -0.06219758520374837, 4.213801391108748, 5.507394037457768, -0.310488259713732, -0.05614154427142712, 6.914605614918611, 5.2859581992078155, -0.3829774142141183, -0.04953703537388402, 9.490159050556638, 5.007043320611547, -0.44982002413274885, -0.042469688627054455, 11.912745930888414, 4.674840124971845, -0.5103368994063947, -0.035029058091642695, 14.156885082907731, 4.294086003296922, -0.5639334415784055, -0.027307519478572413, 16.199587468981022, 3.8700010265739313, -0.6101051102832953, -0.01939915364627895, 18.02058056976475, 3.408219442116292, -0.6484417557795994, -0.011398629051431363},
		'{27.674164915299137, -2.518473327481149, -0.7343556810658288, 0.07050651561734744, 26.267303371140297, -3.10182366472914, -0.673031916650287, 0.07499828955146777, 24.579944291485468, -3.63950419869313, -0.6049442691826482, 0.07854674905513719, 22.6363148619022, -4.126055709312688, -0.5309940973721673, 0.0811266116007131, 20.463203071190655, -4.556702195122791, -0.45213553056660705, 0.08272422960131058, 18.08960476601513, -4.927394718959372, -0.36936354111142766, 0.08333755360923549, 15.546351057643417, -5.234846103754137, -0.2837017436183335, 0.08297596187978151, 12.86572072254922, -5.476556229982458, -0.19619006694069507, 0.08165996051033703, 10.081042334626694, -5.650827799274705, -0.10787244368607801, 0.07942075979238758, 7.226290906312207, -5.756772541325604, -0.019784659468584098, 0.07629973375248308, 4.335683799494449, -5.7943079522396985, 0.06705750012586148, 0.07234777109356638, 1.443280595846728, -5.7641447605759, 0.15166967264396847, 0.06762452686765819, -1.4174085081226995, -5.667765421397324, 0.2331097869118908, 0.06219758520374241, -4.213801391107234, -5.507394037457875, 0.310488259713761, 0.056141544271421234, -6.914605614917137, -5.28595819920792, 0.38297741421414655, 0.04953703537387829, -9.49015905055522, -5.0070433206116505, 0.44982002413277594, 0.04246968862704894, -11.912745930887068, -4.674840124971943, 0.5103368994064205, 0.035029058091637456, -14.156885082906472, -4.294086003297015, 0.5639334415784296, 0.02730751947856751, -16.199587468979864, -3.8700010265740183, 0.6101051102833174, 0.01939915364627442, -18.020580569763702, -3.408219442116372, 0.6484417557796194, 0.011398629051427259},
		'{72.51131969922037, -3.8625231707022207, 0.929323822626333, -0.06994708325861936, 70.5421336889876, -4.011603326911038, 0.9256587549077067, -0.07637552839346037, 68.50214369362797, -4.145796515909857, 0.9201421065661662, -0.082371192286889, 66.39871179008813, -4.265431518949687, 0.9128628483284804, -0.08793909836754918, 64.23903113887704, -4.370854958184794, 0.903910065718909, -0.0930849871807982, 62.03011743793533, -4.462429804040693, 0.8933727614134688, -0.09781527412782093, 59.77880111623674, -4.54053390928278, 0.8813396659957791, -0.10213700750176719, 57.49172025324865, -4.605558571848607, 0.8678990571746913, -0.10605782689940811, 55.1753142093852, -4.657907128358656, 0.8531385875030785, -0.10958592208272783, 52.83581795166512, -4.697993580074422, 0.8371451206171207, -0.11272999236079786, 50.479257057937836, -4.7262412529287605, 0.8200045759961625, -0.11549920655822801, 48.11144338226526, -4.743081493112122, 0.8018017822247844, -0.11790316363245998, 45.7379713633386, -4.748952399559536, 0.7826203387210673, -0.11995185399817505, 43.36421495717219, -4.7442975945474615, 0.7625424858782165, -0.1216556216131318, 40.99532517474419, -4.729565033476708, 0.7416489835506792, -0.12302512687584188, 38.63622820474926, -4.7052058547881135, 0.7200189978007006, -0.12407131038163734, 36.29162410118614, -4.67167327083134, 0.6977299958068675, -0.1248053575798879, 33.96598601512404, -4.6294215003843755, 0.6748576488226227, -0.12523866437139655, 31.66355994967266, -4.578904743402131, 0.6514757430599522, -0.1253828036813429, 29.388365016920893, -4.520576198457048, 0.6276560983614967, -0.12524949303956054},
		'{-72.51131969922082, 3.8625231707022434, -0.9293238226263425, 0.06994708325862117, -70.54213368898823, 4.011603326911068, -0.925658754907719, 0.07637552839346275, -68.50214369362877, 4.145796515909895, -0.9201421065661813, 0.08237119228689191, -66.39871179008907, 4.265431518949732, -0.912862848328498, 0.08793909836755259, -64.2390311388781, 4.370854958184845, -0.903910065718929, 0.09308498718080209, -62.03011743793654, 4.46242980404075, -0.8933727614134911, 0.09781527412782526, -59.778801116238064, 4.540533909282843, -0.8813396659958035, 0.10213700750177193, -57.491720253250094, 4.605558571848675, -0.8678990571747176, 0.10605782689941325, -55.175314209386755, 4.65790712835873, -0.8531385875031068, 0.10958592208273332, -52.83581795166677, 4.697993580074499, -0.8371451206171505, 0.1127299923608037, -50.47925705793958, 4.726241252928842, -0.8200045759961939, 0.11549920655823415, -48.11144338226708, 4.743081493112207, -0.8018017822248172, 0.11790316363246642, -45.737971363340506, 4.7489523995596254, -0.7826203387211014, 0.11995185399818173, -43.36421495717416, 4.744297594547554, -0.7625424858782519, 0.12165562161313871, -40.995325174746235, 4.729565033476804, -0.7416489835507156, 0.12302512687584899, -38.63622820475136, 4.705205854788212, -0.7200189978007379, 0.12407131038164465, -36.29162410118829, 4.671673270831441, -0.6977299958069055, 0.12480535757989536, -33.96598601512623, 4.6294215003844785, -0.6748576488226614, 0.12523866437140418, -31.663559949674887, 4.5789047434022345, -0.6514757430599915, 0.12538280368135063, -29.388365016923153, 4.520576198457154, -0.6276560983615366, 0.12524949303956834}};
	localparam real Fbr[0:3][0:79] = '{
		'{-9.517403442589092, 5.803958733344014, 0.4775028600506327, -0.051475557707039, -12.334175399393775, 5.453185696094708, 0.5490632879926326, -0.04322707994592666, -14.96102263415146, 5.045163100567296, 0.6130702424751429, -0.03461632419982426, -17.37071831975333, 4.585572275315287, 0.6689092796911043, -0.025749026363305512, -19.53900499187631, 4.080596352735773, 0.7160707871752784, -0.01673212178091013, -21.444825625147537, 3.5368402976503113, 0.7541541277356487, -0.007672487370335698, -23.070513795269598, 2.9612473918572286, 0.7828704526032709, 0.0013242945205483789, -24.401941410865636, 2.3610132006917723, 0.8020441735158046, 0.010155136578104976, -25.428623015324696, 1.7434980596004206, 0.8116130991452264, 0.018720598010421204, -26.143776178374335, 1.1161391184899858, 0.8116272566501304, 0.02692597454909598, -26.544338013417295, 0.486362969358328, 0.802246434005084, 0.03468231537764404, -26.630938363918823, -0.1385001412055984, 0.7837364929699213, 0.04190735643865942, -26.407830694600133, -0.7512995481769507, 0.7564645159572013, 0.048526360716390216, -25.882782195429897, -1.345143932141644, 0.7208928624949469, 0.05447285732557144, -25.066925053280514, -1.913476746075026, 0.677572222336209, 0.05968927254545548, -23.974571262882375, -2.4501465043811197, 0.6271337624237217, 0.06412744730359313, -22.622993731046726, -2.949471206591621, 0.5702804737794054, 0.06774903702028089, -21.03217677218664, -3.406296248196691, 0.5077778318738266, 0.0705257911547416, -19.224539395604726, -3.8160452573072905, 0.4404438900763632, 0.07243971123109369, -17.224635043031086, -4.174763387130108, 0.36913893034683815, 0.0734830875492399},
		'{-9.51740344258746, 5.803958733344131, 0.47750286005066395, -0.05147555770703265, -12.334175399392215, 5.45318569609482, 0.5490632879926624, -0.043227079945920587, -14.961022634149993, 5.045163100567405, 0.613070242475171, -0.03461632419981855, -17.37071831975197, 4.585572275315388, 0.6689092796911302, -0.0257490263633002, -19.53900499187507, 4.080596352735866, 0.716070787175302, -0.016732121780905287, -21.444825625146432, 3.5368402976503965, 0.7541541277356698, -0.0076724873703313615, -23.07051379526864, 2.961247391857304, 0.7828704526032892, 0.0013242945205521675, -24.401941410864822, 2.361013200691838, 0.8020441735158201, 0.010155136578108175, -25.428623015324046, 1.743498059600476, 0.8116130991452388, 0.018720598010423785, -26.143776178373848, 1.1161391184900298, 0.8116272566501396, 0.026925974549097925, -26.544338013416983, 0.4863629693583609, 0.8022464340050901, 0.03468231537764534, -26.63093836391867, -0.1385001412055773, 0.7837364929699241, 0.041907356438660066, -26.407830694600147, -0.7512995481769416, 0.7564645159572009, 0.04852636071639022, -25.882782195430078, -1.3451439321416463, 0.7208928624949434, 0.054472857325570806, -25.06692505328085, -1.9134767460750393, 0.6775722223362024, 0.05968927254545422, -23.974571262882865, -2.450146504381144, 0.6271337624237122, 0.0641274473035913, -22.62299373104736, -2.949471206591656, 0.5702804737793931, 0.06774903702027849, -21.032176772187412, -3.406296248196736, 0.507777831873812, 0.07052579115473867, -19.224539395605618, -3.8160452573073442, 0.44044389007634605, 0.07243971123109028, -17.224635043032087, -4.17476338713017, 0.3691389303468188, 0.07348308754923608},
		'{9.313313592773765, -5.688953814066472, -0.40599510904134345, -0.19382811981932202, 12.087015729293103, -5.405857783345071, -0.3589502986526131, -0.18671439091601966, 14.719161330735629, -5.1228350901578645, -0.31308546179083796, -0.17949236217734052, 17.209940666047885, -4.8404954274546945, -0.2684508079689891, -0.17218217464535937, 19.559842146665797, -4.559421645725951, -0.22509179460033948, -0.16480332234289366, 21.769638866145826, -4.280169607798952, -0.18304922627424028, -0.1573746369854663, 23.840375083421378, -4.003268108103177, -0.14235935997530536, -0.14991427476315658, 25.77335268129348, -3.7292188538971804, -0.10305401577095727, -0.14243970513484921, 27.570117630503294, -3.4584965059201647, -0.0651606925002054, -0.13496770157542248, 29.23244648845956, -3.191548775908135, -0.0287026880051382, -0.1275143342146665, 30.762332960409537, -2.9287965783978374, 0.006300776544155451, -0.12009496430516839, 32.16197454955081, -2.6706342342314704, 0.039834428670685595, -0.11272424045505701, 33.43375932128638, -2.417429723170744, 0.07188681338676661, -0.10541609656034238, 34.58025280553011, -2.169524983030432, 0.10245015918354083, -0.09818375137062299, 35.60418505967578, -1.927236252748512, 0.13152024162071368, -0.09103970962115071, 36.508437913554964, -1.6908544568223671, 0.15909624491166258, -0.0839957646636417, 37.2960324164273, -1.4606456285578837, 0.18518062188698006, -0.07706300252778789, 37.9701165047758, -1.2368513696004657, 0.2097789527070889, -0.07025180734515825, 38.53395290842061, -1.0196893432437162, 0.23289980268185642, -0.06357186806706984, 38.990907311220546, -0.8093537990426116, 0.2545545795421773, -0.05703218640805522},
		'{9.313313592769488, -5.688953814066671, -0.40599510904141745, -0.1938281198193366, 12.08701572928894, -5.405857783345265, -0.35895029865268496, -0.18671439091603384, 14.71916133073158, -5.122835090158053, -0.31308546179090785, -0.1794923621773543, 17.209940666043956, -4.8404954274548775, -0.2684508079690569, -0.17218217464537272, 19.559842146661993, -4.559421645726127, -0.22509179460040502, -0.1648033223429066, 21.769638866142145, -4.280169607799123, -0.18304922627430356, -0.15737463698547874, 23.84037508341783, -4.0032681081033425, -0.14235935997536636, -0.14991427476316863, 25.773352681290067, -3.729218853897339, -0.10305401577101594, -0.14243970513486076, 27.570117630500015, -3.4584965059203165, -0.06516069250026163, -0.13496770157543359, 29.232446488456414, -3.191548775908281, -0.0287026880051921, -0.12751433421467714, 30.76233296040653, -2.9287965783979777, 0.0063007765441039365, -0.12009496430517856, 32.161974549547935, -2.6706342342316036, 0.039834428670636524, -0.1127242404550667, 33.43375932128365, -2.41742972317087, 0.07188681338671998, -0.10541609656035161, 34.580252805527515, -2.169524983030552, 0.10245015918349654, -0.09818375137063172, 35.60418505967332, -1.9272362527486258, 0.13152024162067183, -0.09103970962115898, 36.50843791355265, -1.6908544568224744, 0.1590962449116232, -0.0839957646636495, 37.29603241642513, -1.4606456285579843, 0.1851806218869431, -0.0770630025277952, 37.97011650477375, -1.23685136960056, 0.2097789527070543, -0.0702518073451651, 38.5339529084187, -1.0196893432438041, 0.23289980268182417, -0.06357186806707624, 38.99090731121877, -0.8093537990426936, 0.25455457954214733, -0.05703218640806115}};
	localparam real Fbi[0:3][0:79] = '{
		'{27.674164915298654, 2.5184733274811264, -0.7343556810658382, -0.07050651561734925, 26.267303371139647, 3.101823664729105, -0.6730319166502996, -0.07499828955147023, 24.57994429148466, 3.639504198693084, -0.6049442691826638, -0.07854674905514027, 22.636314861901248, 4.12605570931263, -0.5309940973721856, -0.08112661160071676, 20.463203071189568, 4.556702195122724, -0.4521355305666279, -0.08272422960131473, 18.089604766013927, 4.927394718959295, -0.3693635411114507, -0.0833375536092401, 15.546351057642116, 5.234846103754052, -0.2837017436183584, -0.08297596187978651, 12.865720722547834, 5.476556229982367, -0.1961900669407216, -0.08165996051034236, 10.081042334625243, 5.650827799274608, -0.10787244368610588, -0.07942075979239319, 7.226290906310707, 5.756772541325502, -0.01978465946861291, -0.07629973375248889, 4.335683799492918, 5.794307952239594, 0.06705750012583211, -0.0723477710935723, 1.4432805958451844, 5.764144760575793, 0.15166967264393882, -0.06762452686766418, -1.4174085081242387, 5.667765421397218, 0.2331097869118613, -0.06219758520374837, -4.213801391108748, 5.507394037457768, 0.310488259713732, -0.05614154427142712, -6.914605614918611, 5.2859581992078155, 0.3829774142141183, -0.04953703537388402, -9.490159050556638, 5.007043320611547, 0.44982002413274885, -0.042469688627054455, -11.912745930888414, 4.674840124971845, 0.5103368994063947, -0.035029058091642695, -14.156885082907731, 4.294086003296922, 0.5639334415784055, -0.027307519478572413, -16.199587468981022, 3.8700010265739313, 0.6101051102832953, -0.01939915364627895, -18.02058056976475, 3.408219442116292, 0.6484417557795994, -0.011398629051431363},
		'{-27.674164915299137, -2.518473327481149, 0.7343556810658288, 0.07050651561734744, -26.267303371140297, -3.10182366472914, 0.673031916650287, 0.07499828955146777, -24.579944291485468, -3.63950419869313, 0.6049442691826482, 0.07854674905513719, -22.6363148619022, -4.126055709312688, 0.5309940973721673, 0.0811266116007131, -20.463203071190655, -4.556702195122791, 0.45213553056660705, 0.08272422960131058, -18.08960476601513, -4.927394718959372, 0.36936354111142766, 0.08333755360923549, -15.546351057643417, -5.234846103754137, 0.2837017436183335, 0.08297596187978151, -12.86572072254922, -5.476556229982458, 0.19619006694069507, 0.08165996051033703, -10.081042334626694, -5.650827799274705, 0.10787244368607801, 0.07942075979238758, -7.226290906312207, -5.756772541325604, 0.019784659468584098, 0.07629973375248308, -4.335683799494449, -5.7943079522396985, -0.06705750012586148, 0.07234777109356638, -1.443280595846728, -5.7641447605759, -0.15166967264396847, 0.06762452686765819, 1.4174085081226995, -5.667765421397324, -0.2331097869118908, 0.06219758520374241, 4.213801391107234, -5.507394037457875, -0.310488259713761, 0.056141544271421234, 6.914605614917137, -5.28595819920792, -0.38297741421414655, 0.04953703537387829, 9.49015905055522, -5.0070433206116505, -0.44982002413277594, 0.04246968862704894, 11.912745930887068, -4.674840124971943, -0.5103368994064205, 0.035029058091637456, 14.156885082906472, -4.294086003297015, -0.5639334415784296, 0.02730751947856751, 16.199587468979864, -3.8700010265740183, -0.6101051102833174, 0.01939915364627442, 18.020580569763702, -3.408219442116372, -0.6484417557796194, 0.011398629051427259},
		'{-72.51131969922037, -3.8625231707022207, -0.929323822626333, -0.06994708325861936, -70.5421336889876, -4.011603326911038, -0.9256587549077067, -0.07637552839346037, -68.50214369362797, -4.145796515909857, -0.9201421065661662, -0.082371192286889, -66.39871179008813, -4.265431518949687, -0.9128628483284804, -0.08793909836754918, -64.23903113887704, -4.370854958184794, -0.903910065718909, -0.0930849871807982, -62.03011743793533, -4.462429804040693, -0.8933727614134688, -0.09781527412782093, -59.77880111623674, -4.54053390928278, -0.8813396659957791, -0.10213700750176719, -57.49172025324865, -4.605558571848607, -0.8678990571746913, -0.10605782689940811, -55.1753142093852, -4.657907128358656, -0.8531385875030785, -0.10958592208272783, -52.83581795166512, -4.697993580074422, -0.8371451206171207, -0.11272999236079786, -50.479257057937836, -4.7262412529287605, -0.8200045759961625, -0.11549920655822801, -48.11144338226526, -4.743081493112122, -0.8018017822247844, -0.11790316363245998, -45.7379713633386, -4.748952399559536, -0.7826203387210673, -0.11995185399817505, -43.36421495717219, -4.7442975945474615, -0.7625424858782165, -0.1216556216131318, -40.99532517474419, -4.729565033476708, -0.7416489835506792, -0.12302512687584188, -38.63622820474926, -4.7052058547881135, -0.7200189978007006, -0.12407131038163734, -36.29162410118614, -4.67167327083134, -0.6977299958068675, -0.1248053575798879, -33.96598601512404, -4.6294215003843755, -0.6748576488226227, -0.12523866437139655, -31.66355994967266, -4.578904743402131, -0.6514757430599522, -0.1253828036813429, -29.388365016920893, -4.520576198457048, -0.6276560983614967, -0.12524949303956054},
		'{72.51131969922082, 3.8625231707022434, 0.9293238226263425, 0.06994708325862117, 70.54213368898823, 4.011603326911068, 0.925658754907719, 0.07637552839346275, 68.50214369362877, 4.145796515909895, 0.9201421065661813, 0.08237119228689191, 66.39871179008907, 4.265431518949732, 0.912862848328498, 0.08793909836755259, 64.2390311388781, 4.370854958184845, 0.903910065718929, 0.09308498718080209, 62.03011743793654, 4.46242980404075, 0.8933727614134911, 0.09781527412782526, 59.778801116238064, 4.540533909282843, 0.8813396659958035, 0.10213700750177193, 57.491720253250094, 4.605558571848675, 0.8678990571747176, 0.10605782689941325, 55.175314209386755, 4.65790712835873, 0.8531385875031068, 0.10958592208273332, 52.83581795166677, 4.697993580074499, 0.8371451206171505, 0.1127299923608037, 50.47925705793958, 4.726241252928842, 0.8200045759961939, 0.11549920655823415, 48.11144338226708, 4.743081493112207, 0.8018017822248172, 0.11790316363246642, 45.737971363340506, 4.7489523995596254, 0.7826203387211014, 0.11995185399818173, 43.36421495717416, 4.744297594547554, 0.7625424858782519, 0.12165562161313871, 40.995325174746235, 4.729565033476804, 0.7416489835507156, 0.12302512687584899, 38.63622820475136, 4.705205854788212, 0.7200189978007379, 0.12407131038164465, 36.29162410118829, 4.671673270831441, 0.6977299958069055, 0.12480535757989536, 33.96598601512623, 4.6294215003844785, 0.6748576488226614, 0.12523866437140418, 31.663559949674887, 4.5789047434022345, 0.6514757430599915, 0.12538280368135063, 29.388365016923153, 4.520576198457154, 0.6276560983615366, 0.12524949303956834}};
endpackage
`endif
