`ifndef COEFFICIENTS_FX_SV_
`define COEFFICIENTS_FX_SV_

package Coefficients_Fx;

	localparam N = 4;
	localparam COEFF_BIAS = 48;
	localparam logic signed[63:0] Lfr[0:3] = {64'd272579065432618, 64'd272579065432618, 64'd264866559397522, 64'd264866559397522};

	localparam logic signed[63:0] Lfi[0:3] = {64'd33142944436156, - 64'd33142944436156, 64'd12931747597259, - 64'd12931747597259};

	localparam logic signed[63:0] Lbr[0:3] = {64'd272579065432618, 64'd272579065432618, 64'd264866559397522, 64'd264866559397522};

	localparam logic signed[63:0] Lbi[0:3] = {64'd33142944436156, - 64'd33142944436156, 64'd12931747597259, - 64'd12931747597259};

	localparam logic signed[63:0] Wfr[0:3] = {- 64'd142796336093, - 64'd142796336093, 64'd41600396254, 64'd41600396254};

	localparam logic signed[63:0] Wfi[0:3] = {- 64'd10038173912, 64'd10038173912, 64'd83875608999, - 64'd83875608999};

	localparam logic signed[63:0] Wbr[0:3] = {64'd142796336093, 64'd142796336093, - 64'd41600396254, - 64'd41600396254};

	localparam logic signed[63:0] Wbi[0:3] = {64'd10038173912, - 64'd10038173912, - 64'd83875608999, 64'd83875608999};

	localparam logic signed[63:0] Ffr[0:3][0:79] = '{
		'{- 64'd3416995017050702, - 64'd790736473211221, 64'd228205129574949, - 64'd5800094494514, - 64'd3776115705624860, - 64'd645233420583674, 64'd229585273724347, - 64'd10349661644996, - 64'd4061748819895167, - 64'd497174553008282, 64'd227486298533109, - 64'd14525445513296, - 64'd4273201735636153, - 64'd348884077258512, 64'd222107603032668, - 64'd18283451076243, - 64'd4410917876795718, - 64'd202577276583765, 64'd213687693587887, - 64'd21588019856460, - 64'd4476415201422712, - 64'd60332850299622, 64'd202498748224028, - 64'd24411956886811, - 64'd4472211690427369, 64'd75931379265017, 64'd188840943274486, - 64'd26736525740924, - 64'd4401739575017963, 64'd204479194187039, 64'd173036638164860, - 64'd28551318082134, - 64'd4269250122116482, 64'd323773007040548, 64'd155424511625192, - 64'd29854005736309, - 64'd4079710849439797, 64'd432487111540906, 64'd136353738833879, - 64'd30649984653062, - 64'd3838697063964515, 64'd529517143320681, 64'd116178294061222, - 64'd30951921274023, - 64'd3552279610313324, 64'd613985793443917, 64'd95251457426747, - 64'd30779212768861, - 64'd3226910680727266, 64'd685244870901960, 64'd73920597549936, - 64'd30157373325874, - 64'd2869309477579148, 64'd742873859947327, 64'd52522294303071, - 64'd29117359193852, - 64'd2486349434989546, 64'd786675163168762, 64'd31377857715622, - 64'd27694845468458, - 64'd2084948600428164, 64'd816666261242094, 64'd10789290481732, - 64'd25929467705413, - 64'd1671964652819259, 64'd833069054955107, - 64'd8964267365161, - 64'd23864041333108, - 64'd1254095893372400, 64'd836296684144756, - 64'd27629582077513, - 64'd21543771540048, - 64'd837789391984547, 64'd826938141441906, - 64'd44981837618987, - 64'd19015465841321, - 64'd429157308518182, 64'd805741016126249, - 64'd60826603291541, - 64'd16326760898421},
		'{- 64'd3416995017050815, - 64'd790736473211198, 64'd228205129574948, - 64'd5800094494514, - 64'd3776115705624978, - 64'd645233420583651, 64'd229585273724345, - 64'd10349661644995, - 64'd4061748819895286, - 64'd497174553008260, 64'd227486298533108, - 64'd14525445513296, - 64'd4273201735636272, - 64'd348884077258492, 64'd222107603032667, - 64'd18283451076242, - 64'd4410917876795836, - 64'd202577276583746, 64'd213687693587886, - 64'd21588019856460, - 64'd4476415201422826, - 64'd60332850299605, 64'd202498748224027, - 64'd24411956886811, - 64'd4472211690427478, 64'd75931379265032, 64'd188840943274485, - 64'd26736525740924, - 64'd4401739575018065, 64'd204479194187053, 64'd173036638164858, - 64'd28551318082134, - 64'd4269250122116577, 64'd323773007040559, 64'd155424511625190, - 64'd29854005736309, - 64'd4079710849439883, 64'd432487111540915, 64'd136353738833878, - 64'd30649984653062, - 64'd3838697063964592, 64'd529517143320688, 64'd116178294061221, - 64'd30951921274023, - 64'd3552279610313391, 64'd613985793443922, 64'd95251457426746, - 64'd30779212768861, - 64'd3226910680727322, 64'd685244870901963, 64'd73920597549935, - 64'd30157373325874, - 64'd2869309477579193, 64'd742873859947328, 64'd52522294303070, - 64'd29117359193852, - 64'd2486349434989580, 64'd786675163168761, 64'd31377857715621, - 64'd27694845468458, - 64'd2084948600428186, 64'd816666261242091, 64'd10789290481732, - 64'd25929467705413, - 64'd1671964652819271, 64'd833069054955102, - 64'd8964267365162, - 64'd23864041333108, - 64'd1254095893372402, 64'd836296684144750, - 64'd27629582077514, - 64'd21543771540049, - 64'd837789391984538, 64'd826938141441898, - 64'd44981837618987, - 64'd19015465841322, - 64'd429157308518163, 64'd805741016126240, - 64'd60826603291541, - 64'd16326760898421},
		'{64'd3275922003959216, 64'd760659500307872, - 64'd202576595739189, 64'd72238367289273, 64'd3624719872900220, 64'd636449918759182, - 64'd175271156122064, 64'd65744873177707, 64'd3914036119240986, 64'd522644442827493, - 64'd150055154649368, 64'd59613695258635, 64'd4148939572491594, 64'd418709905349560, - 64'd126834717817234, 64'd53838390361862, 64'd4334233530640439, 64'd324117875028896, - 64'd105515365308010, 64'd48411249485237, 64'd4474458748962082, 64'd238347079200576, - 64'd86002606571427, 64'd43323483207658, 64'd4573897561054708, 64'd160885514201279, - 64'd68202470396773, 64'd38565392300456, 64'd4636578981778483, 64'd91232266661397, - 64'd52021972047535, 64'd34126524246988, 64'd4666284653174622, 64'd28899068031350, - 64'd37369522365210, 64'd29995816379323, 64'd4666555505347799, - 64'd26588396362110, - 64'd24155283078135, 64'd26161726335999, 64'd4640699014687624, - 64'd75689403455150, - 64'd12291472375824, 64'd22612350536644, 64'd4591796951687465, - 64'd118847314527012, - 64'd1692624630987, 64'd19335531358022, 64'd4522713519992917, - 64'd156488884979320, 64'd7724192028627, 64'd16318953682290, 64'd4436103797182666, - 64'd189023744573788, 64'd16039196776865, 64'd13550231472305, 64'd4334422396158091, - 64'd216844031872483, 64'd23329752432474, 64'd11016985010939, 64'd4219932273904040, - 64'd240324167589901, 64'd29670253925608, 64'd8706909422000, 64'd4094713621792180, - 64'd259820752508214, 64'd35132045900064, 64'd6607835069660, 64'd3960672778542676, - 64'd275672576523485, 64'd39783366636658, 64'd4707780411615, 64'd3819551113452787, - 64'd288200726279196, 64'd43689315652394, 64'd2994997858749, 64'd3672933833557044, - 64'd297708779702204, 64'd46911842495046, 64'd1458013171010},
		'{64'd3275922003959475, 64'd760659500307814, - 64'd202576595739187, 64'd72238367289273, 64'd3624719872900466, 64'd636449918759128, - 64'd175271156122062, 64'd65744873177707, 64'd3914036119241220, 64'd522644442827442, - 64'd150055154649366, 64'd59613695258634, 64'd4148939572491815, 64'd418709905349512, - 64'd126834717817232, 64'd53838390361861, 64'd4334233530640648, 64'd324117875028852, - 64'd105515365308008, 64'd48411249485236, 64'd4474458748962279, 64'd238347079200534, - 64'd86002606571426, 64'd43323483207658, 64'd4573897561054892, 64'd160885514201241, - 64'd68202470396772, 64'd38565392300455, 64'd4636578981778655, 64'd91232266661362, - 64'd52021972047533, 64'd34126524246988, 64'd4666284653174782, 64'd28899068031317, - 64'd37369522365208, 64'd29995816379323, 64'd4666555505347949, - 64'd26588396362141, - 64'd24155283078133, 64'd26161726335998, 64'd4640699014687764, - 64'd75689403455178, - 64'd12291472375823, 64'd22612350536644, 64'd4591796951687594, - 64'd118847314527037, - 64'd1692624630986, 64'd19335531358021, 64'd4522713519993036, - 64'd156488884979343, 64'd7724192028628, 64'd16318953682290, 64'd4436103797182776, - 64'd189023744573809, 64'd16039196776866, 64'd13550231472305, 64'd4334422396158192, - 64'd216844031872502, 64'd23329752432475, 64'd11016985010939, 64'd4219932273904134, - 64'd240324167589918, 64'd29670253925609, 64'd8706909422000, 64'd4094713621792266, - 64'd259820752508229, 64'd35132045900065, 64'd6607835069659, 64'd3960672778542754, - 64'd275672576523500, 64'd39783366636659, 64'd4707780411615, 64'd3819551113452858, - 64'd288200726279208, 64'd43689315652395, 64'd2994997858748, 64'd3672933833557108, - 64'd297708779702215, 64'd46911842495047, 64'd1458013171010}};

	localparam logic signed[63:0] Ffi[0:3][0:79] = '{
		'{64'd3967081808774704, - 64'd1023480183090411, - 64'd72973861234924, 64'd40195174460707, 64'd3439361421235583, - 64'd1084240632532636, - 64'd43796990805152, 64'd38241875017222, 64'd2886033914497596, - 64'd1125948165731119, - 64'd15379736069659, 64'd35814609204551, 64'd2316561562200497, - 64'd1148904002427228, 64'd11892253112228, 64'd32972368559049, 64'd1740189141063770, - 64'd1153673511711328, 64'd37668993916565, 64'd29777460510886, 64'd1165817038085718, - 64'd1141065038220589, 64'd61639648098001, 64'd26294421979944, 64'd601885611263630, - 64'd1112106140585773, 64'd83535249590230, 64'd22588952357362, 64'd56271978554240, - 64'd1068017720409403, 64'd103130677879204, 64'd18726880794959, - 64'd463799831723903, - 64'd1010186528288342, 64'd120245884282124, 64'd14773181493349, - 64'd951834679556170, - 64'd940136533995375, 64'd134746389024622, 64'd10791049304289, - 64'd1402127613652993, - 64'd859499641266716, 64'd146543076981889, 64'd6841046470907, - 64'd1809810463431250, - 64'd769986214155986, 64'd155591329026457, 64'd2980329748836, - 64'd2170883741138742, - 64'd673355862140346, 64'd161889534014421, - 64'd738034490298, - 64'd2482234090146021, - 64'd571388905698901, 64'd165477033470502, - 64'd4265661246813, - 64'd2741637718850605, - 64'd465858913581007, 64'd166431556947436, - 64'd7559339728395, - 64'd2947750446693363, - 64'd358506668139424, 64'd164866210802551, - 64'd10581425453121, - 64'd3100085157486249, - 64'd251015876648266, 64'd160926086738719, - 64'd13300130662146, - 64'd3198977603974878, - 64'd144990905204435, 64'd154784558900808, - 64'd15689713641879, - 64'd3245541635063636, - 64'd41936768376526, 64'd146639339622087, - 64'd17730569029005, - 64'd3241615022545980, 64'd56758437035178, 64'd136708364113511, - 64'd19409222543207},
		'{- 64'd3967081808774766, 64'd1023480183090412, 64'd72973861234923, - 64'd40195174460707, - 64'd3439361421235630, 64'd1084240632532635, 64'd43796990805150, - 64'd38241875017222, - 64'd2886033914497626, 64'd1125948165731114, 64'd15379736069658, - 64'd35814609204551, - 64'd2316561562200513, 64'd1148904002427221, - 64'd11892253112229, - 64'd32972368559049, - 64'd1740189141063773, 64'd1153673511711319, - 64'd37668993916565, - 64'd29777460510887, - 64'd1165817038085706, 64'd1141065038220578, - 64'd61639648098002, - 64'd26294421979944, - 64'd601885611263606, 64'd1112106140585761, - 64'd83535249590230, - 64'd22588952357362, - 64'd56271978554203, 64'd1068017720409389, - 64'd103130677879204, - 64'd18726880794959, 64'd463799831723951, 64'd1010186528288326, - 64'd120245884282124, - 64'd14773181493349, 64'd951834679556227, 64'd940136533995359, - 64'd134746389024622, - 64'd10791049304289, 64'd1402127613653059, 64'd859499641266700, - 64'd146543076981888, - 64'd6841046470907, 64'd1809810463431322, 64'd769986214155970, - 64'd155591329026456, - 64'd2980329748836, 64'd2170883741138821, 64'd673355862140328, - 64'd161889534014420, 64'd738034490298, 64'd2482234090146103, 64'd571388905698884, - 64'd165477033470501, 64'd4265661246813, 64'd2741637718850690, 64'd465858913580991, - 64'd166431556947434, 64'd7559339728395, 64'd2947750446693449, 64'd358506668139408, - 64'd164866210802549, 64'd10581425453120, 64'd3100085157486335, 64'd251015876648252, - 64'd160926086738718, 64'd13300130662146, 64'd3198977603974963, 64'd144990905204422, - 64'd154784558900806, 64'd15689713641879, 64'd3245541635063718, 64'd41936768376513, - 64'd146639339622086, 64'd17730569029005, 64'd3241615022546059, - 64'd56758437035189, - 64'd136708364113510, 64'd19409222543207},
		'{- 64'd11799314100150670, 64'd1726645102791665, - 64'd334163755354307, 64'd48561971159818, - 64'd10952591127214628, 64'd1659711317154405, - 64'd323753374549305, 64'd49015407026636, - 64'd10139804252581744, 64'd1591020420745462, - 64'd312702769499617, 64'd49143758653124, - 64'd9361683830509244, 64'd1521154085508429, - 64'd301145711237301, 64'd48982853438203, - 64'd8618684244533847, 64'd1450635166671628, - 64'd289203764829884, 64'd48566108769607, - 64'd7911012390371385, 64'd1379931390804498, - 64'd276986981713980, 64'd47924616070612, - 64'd7238654340870150, 64'd1309458937568988, - 64'd264594578586406, 64'd47087228405991, - 64'd6601400248267951, 64'd1239585907086178, - 64'd252115600567391, 64'd46080650757144, - 64'd5998867542649463, 64'd1170635666386360, - 64'd239629566695339, 64'd44929532161494, - 64'd5430522488407580, 64'd1102890069821280, - 64'd227207096129585, 64'd43656558991310, - 64'd4895700162747228, 64'd1036592549597817, - 64'd214910513727958, 64'd42282548722202, - 64'd4393622921895572, 64'd971951073750469, - 64'd202794433931221, 64'd40826543611873, - 64'd3923417421757894, 64'd909140969912908, - 64'd190906322127786, 64'd39305903775323, - 64'd3484130260339856, 64'd848307614183701, - 64'd179287032890993, 64'd37736399203861, - 64'd3074742309396342, 64'd789568985214973, - 64'd167971324678882, 64'd36132300332036, - 64'd2694181802513566, 64'd733018084392030, - 64'd156988350764125, 64'd34506466809278, - 64'd2341336246230446, 64'd678725223623238, - 64'd146362126320812, 64'd32870434181603, - 64'd2015063219899441, 64'd626740182829036, - 64'd136111971736398, 64'd31234498233591, - 64'd1714200128815726, 64'd577094239712797, - 64'd126252932342361, 64'd29607796781994, - 64'd1437572973743111, 64'd529802074820183, - 64'd116796174867260, 64'd27998388750033},
		'{64'd11799314100150724, - 64'd1726645102791664, 64'd334163755354309, - 64'd48561971159818, 64'd10952591127214666, - 64'd1659711317154402, 64'd323753374549306, - 64'd49015407026636, 64'd10139804252581770, - 64'd1591020420745457, 64'd312702769499617, - 64'd49143758653124, 64'd9361683830509258, - 64'd1521154085508422, 64'd301145711237302, - 64'd48982853438203, 64'd8618684244533850, - 64'd1450635166671619, 64'd289203764829885, - 64'd48566108769607, 64'd7911012390371378, - 64'd1379931390804488, 64'd276986981713981, - 64'd47924616070612, 64'd7238654340870134, - 64'd1309458937568976, 64'd264594578586406, - 64'd47087228405991, 64'd6601400248267928, - 64'd1239585907086164, 64'd252115600567391, - 64'd46080650757144, 64'd5998867542649432, - 64'd1170635666386346, 64'd239629566695339, - 64'd44929532161494, 64'd5430522488407544, - 64'd1102890069821265, 64'd227207096129585, - 64'd43656558991310, 64'd4895700162747188, - 64'd1036592549597802, 64'd214910513727958, - 64'd42282548722202, 64'd4393622921895528, - 64'd971951073750454, 64'd202794433931221, - 64'd40826543611872, 64'd3923417421757846, - 64'd909140969912892, 64'd190906322127786, - 64'd39305903775323, 64'd3484130260339806, - 64'd848307614183685, 64'd179287032890993, - 64'd37736399203861, 64'd3074742309396289, - 64'd789568985214957, 64'd167971324678882, - 64'd36132300332036, 64'd2694181802513512, - 64'd733018084392014, 64'd156988350764125, - 64'd34506466809278, 64'd2341336246230391, - 64'd678725223623223, 64'd146362126320812, - 64'd32870434181603, 64'd2015063219899384, - 64'd626740182829020, 64'd136111971736398, - 64'd31234498233591, 64'd1714200128815670, - 64'd577094239712781, 64'd126252932342361, - 64'd29607796781994, 64'd1437572973743055, - 64'd529802074820168, 64'd116796174867260, - 64'd27998388750033}};

	localparam logic signed[63:0] Fbr[0:3][0:79] = '{
		'{64'd3416995017050702, - 64'd790736473211221, - 64'd228205129574949, - 64'd5800094494514, 64'd3776115705624860, - 64'd645233420583674, - 64'd229585273724347, - 64'd10349661644996, 64'd4061748819895167, - 64'd497174553008282, - 64'd227486298533109, - 64'd14525445513296, 64'd4273201735636153, - 64'd348884077258512, - 64'd222107603032668, - 64'd18283451076243, 64'd4410917876795718, - 64'd202577276583765, - 64'd213687693587887, - 64'd21588019856460, 64'd4476415201422712, - 64'd60332850299622, - 64'd202498748224028, - 64'd24411956886811, 64'd4472211690427369, 64'd75931379265017, - 64'd188840943274486, - 64'd26736525740924, 64'd4401739575017963, 64'd204479194187039, - 64'd173036638164860, - 64'd28551318082134, 64'd4269250122116482, 64'd323773007040548, - 64'd155424511625192, - 64'd29854005736309, 64'd4079710849439797, 64'd432487111540906, - 64'd136353738833879, - 64'd30649984653062, 64'd3838697063964515, 64'd529517143320681, - 64'd116178294061222, - 64'd30951921274023, 64'd3552279610313324, 64'd613985793443917, - 64'd95251457426747, - 64'd30779212768861, 64'd3226910680727266, 64'd685244870901960, - 64'd73920597549936, - 64'd30157373325874, 64'd2869309477579148, 64'd742873859947327, - 64'd52522294303071, - 64'd29117359193852, 64'd2486349434989546, 64'd786675163168762, - 64'd31377857715622, - 64'd27694845468458, 64'd2084948600428164, 64'd816666261242094, - 64'd10789290481732, - 64'd25929467705413, 64'd1671964652819259, 64'd833069054955107, 64'd8964267365161, - 64'd23864041333108, 64'd1254095893372400, 64'd836296684144756, 64'd27629582077513, - 64'd21543771540048, 64'd837789391984547, 64'd826938141441906, 64'd44981837618987, - 64'd19015465841321, 64'd429157308518182, 64'd805741016126249, 64'd60826603291541, - 64'd16326760898421},
		'{64'd3416995017050815, - 64'd790736473211198, - 64'd228205129574948, - 64'd5800094494514, 64'd3776115705624978, - 64'd645233420583651, - 64'd229585273724345, - 64'd10349661644995, 64'd4061748819895286, - 64'd497174553008260, - 64'd227486298533108, - 64'd14525445513296, 64'd4273201735636272, - 64'd348884077258492, - 64'd222107603032667, - 64'd18283451076242, 64'd4410917876795836, - 64'd202577276583746, - 64'd213687693587886, - 64'd21588019856460, 64'd4476415201422826, - 64'd60332850299605, - 64'd202498748224027, - 64'd24411956886811, 64'd4472211690427478, 64'd75931379265032, - 64'd188840943274485, - 64'd26736525740924, 64'd4401739575018065, 64'd204479194187053, - 64'd173036638164858, - 64'd28551318082134, 64'd4269250122116577, 64'd323773007040559, - 64'd155424511625190, - 64'd29854005736309, 64'd4079710849439883, 64'd432487111540915, - 64'd136353738833878, - 64'd30649984653062, 64'd3838697063964592, 64'd529517143320688, - 64'd116178294061221, - 64'd30951921274023, 64'd3552279610313391, 64'd613985793443922, - 64'd95251457426746, - 64'd30779212768861, 64'd3226910680727322, 64'd685244870901963, - 64'd73920597549935, - 64'd30157373325874, 64'd2869309477579193, 64'd742873859947328, - 64'd52522294303070, - 64'd29117359193852, 64'd2486349434989580, 64'd786675163168761, - 64'd31377857715621, - 64'd27694845468458, 64'd2084948600428186, 64'd816666261242091, - 64'd10789290481732, - 64'd25929467705413, 64'd1671964652819271, 64'd833069054955102, 64'd8964267365162, - 64'd23864041333108, 64'd1254095893372402, 64'd836296684144750, 64'd27629582077514, - 64'd21543771540049, 64'd837789391984538, 64'd826938141441898, 64'd44981837618987, - 64'd19015465841322, 64'd429157308518163, 64'd805741016126240, 64'd60826603291541, - 64'd16326760898421},
		'{- 64'd3275922003959216, 64'd760659500307872, 64'd202576595739189, 64'd72238367289273, - 64'd3624719872900220, 64'd636449918759182, 64'd175271156122064, 64'd65744873177707, - 64'd3914036119240986, 64'd522644442827493, 64'd150055154649368, 64'd59613695258635, - 64'd4148939572491594, 64'd418709905349560, 64'd126834717817234, 64'd53838390361862, - 64'd4334233530640439, 64'd324117875028896, 64'd105515365308010, 64'd48411249485237, - 64'd4474458748962082, 64'd238347079200576, 64'd86002606571427, 64'd43323483207658, - 64'd4573897561054708, 64'd160885514201279, 64'd68202470396773, 64'd38565392300456, - 64'd4636578981778483, 64'd91232266661397, 64'd52021972047535, 64'd34126524246988, - 64'd4666284653174622, 64'd28899068031350, 64'd37369522365210, 64'd29995816379323, - 64'd4666555505347799, - 64'd26588396362110, 64'd24155283078135, 64'd26161726335999, - 64'd4640699014687624, - 64'd75689403455150, 64'd12291472375824, 64'd22612350536644, - 64'd4591796951687465, - 64'd118847314527012, 64'd1692624630987, 64'd19335531358022, - 64'd4522713519992917, - 64'd156488884979320, - 64'd7724192028627, 64'd16318953682290, - 64'd4436103797182666, - 64'd189023744573788, - 64'd16039196776865, 64'd13550231472305, - 64'd4334422396158091, - 64'd216844031872483, - 64'd23329752432474, 64'd11016985010939, - 64'd4219932273904040, - 64'd240324167589901, - 64'd29670253925608, 64'd8706909422000, - 64'd4094713621792180, - 64'd259820752508214, - 64'd35132045900064, 64'd6607835069660, - 64'd3960672778542676, - 64'd275672576523485, - 64'd39783366636658, 64'd4707780411615, - 64'd3819551113452787, - 64'd288200726279196, - 64'd43689315652394, 64'd2994997858749, - 64'd3672933833557044, - 64'd297708779702204, - 64'd46911842495046, 64'd1458013171010},
		'{- 64'd3275922003959475, 64'd760659500307814, 64'd202576595739187, 64'd72238367289273, - 64'd3624719872900466, 64'd636449918759128, 64'd175271156122062, 64'd65744873177707, - 64'd3914036119241220, 64'd522644442827442, 64'd150055154649366, 64'd59613695258634, - 64'd4148939572491815, 64'd418709905349512, 64'd126834717817232, 64'd53838390361861, - 64'd4334233530640648, 64'd324117875028852, 64'd105515365308008, 64'd48411249485236, - 64'd4474458748962279, 64'd238347079200534, 64'd86002606571426, 64'd43323483207658, - 64'd4573897561054892, 64'd160885514201241, 64'd68202470396772, 64'd38565392300455, - 64'd4636578981778655, 64'd91232266661362, 64'd52021972047533, 64'd34126524246988, - 64'd4666284653174782, 64'd28899068031317, 64'd37369522365208, 64'd29995816379323, - 64'd4666555505347949, - 64'd26588396362141, 64'd24155283078133, 64'd26161726335998, - 64'd4640699014687764, - 64'd75689403455178, 64'd12291472375823, 64'd22612350536644, - 64'd4591796951687594, - 64'd118847314527037, 64'd1692624630986, 64'd19335531358021, - 64'd4522713519993036, - 64'd156488884979343, - 64'd7724192028628, 64'd16318953682290, - 64'd4436103797182776, - 64'd189023744573809, - 64'd16039196776866, 64'd13550231472305, - 64'd4334422396158192, - 64'd216844031872502, - 64'd23329752432475, 64'd11016985010939, - 64'd4219932273904134, - 64'd240324167589918, - 64'd29670253925609, 64'd8706909422000, - 64'd4094713621792266, - 64'd259820752508229, - 64'd35132045900065, 64'd6607835069659, - 64'd3960672778542754, - 64'd275672576523500, - 64'd39783366636659, 64'd4707780411615, - 64'd3819551113452858, - 64'd288200726279208, - 64'd43689315652395, 64'd2994997858748, - 64'd3672933833557108, - 64'd297708779702215, - 64'd46911842495047, 64'd1458013171010}};

	localparam logic signed[63:0] Fbi[0:3][0:79] = '{
		'{- 64'd3967081808774704, - 64'd1023480183090411, 64'd72973861234924, 64'd40195174460707, - 64'd3439361421235583, - 64'd1084240632532636, 64'd43796990805152, 64'd38241875017222, - 64'd2886033914497596, - 64'd1125948165731119, 64'd15379736069659, 64'd35814609204551, - 64'd2316561562200497, - 64'd1148904002427228, - 64'd11892253112228, 64'd32972368559049, - 64'd1740189141063770, - 64'd1153673511711328, - 64'd37668993916565, 64'd29777460510886, - 64'd1165817038085718, - 64'd1141065038220589, - 64'd61639648098001, 64'd26294421979944, - 64'd601885611263630, - 64'd1112106140585773, - 64'd83535249590230, 64'd22588952357362, - 64'd56271978554240, - 64'd1068017720409403, - 64'd103130677879204, 64'd18726880794959, 64'd463799831723903, - 64'd1010186528288342, - 64'd120245884282124, 64'd14773181493349, 64'd951834679556170, - 64'd940136533995375, - 64'd134746389024622, 64'd10791049304289, 64'd1402127613652993, - 64'd859499641266716, - 64'd146543076981889, 64'd6841046470907, 64'd1809810463431250, - 64'd769986214155986, - 64'd155591329026457, 64'd2980329748836, 64'd2170883741138742, - 64'd673355862140346, - 64'd161889534014421, - 64'd738034490298, 64'd2482234090146021, - 64'd571388905698901, - 64'd165477033470502, - 64'd4265661246813, 64'd2741637718850605, - 64'd465858913581007, - 64'd166431556947436, - 64'd7559339728395, 64'd2947750446693363, - 64'd358506668139424, - 64'd164866210802551, - 64'd10581425453121, 64'd3100085157486249, - 64'd251015876648266, - 64'd160926086738719, - 64'd13300130662146, 64'd3198977603974878, - 64'd144990905204435, - 64'd154784558900808, - 64'd15689713641879, 64'd3245541635063636, - 64'd41936768376526, - 64'd146639339622087, - 64'd17730569029005, 64'd3241615022545980, 64'd56758437035178, - 64'd136708364113511, - 64'd19409222543207},
		'{64'd3967081808774766, 64'd1023480183090412, - 64'd72973861234923, - 64'd40195174460707, 64'd3439361421235630, 64'd1084240632532635, - 64'd43796990805150, - 64'd38241875017222, 64'd2886033914497626, 64'd1125948165731114, - 64'd15379736069658, - 64'd35814609204551, 64'd2316561562200513, 64'd1148904002427221, 64'd11892253112229, - 64'd32972368559049, 64'd1740189141063773, 64'd1153673511711319, 64'd37668993916565, - 64'd29777460510887, 64'd1165817038085706, 64'd1141065038220578, 64'd61639648098002, - 64'd26294421979944, 64'd601885611263606, 64'd1112106140585761, 64'd83535249590230, - 64'd22588952357362, 64'd56271978554203, 64'd1068017720409389, 64'd103130677879204, - 64'd18726880794959, - 64'd463799831723951, 64'd1010186528288326, 64'd120245884282124, - 64'd14773181493349, - 64'd951834679556227, 64'd940136533995359, 64'd134746389024622, - 64'd10791049304289, - 64'd1402127613653059, 64'd859499641266700, 64'd146543076981888, - 64'd6841046470907, - 64'd1809810463431322, 64'd769986214155970, 64'd155591329026456, - 64'd2980329748836, - 64'd2170883741138821, 64'd673355862140328, 64'd161889534014420, 64'd738034490298, - 64'd2482234090146103, 64'd571388905698884, 64'd165477033470501, 64'd4265661246813, - 64'd2741637718850690, 64'd465858913580991, 64'd166431556947434, 64'd7559339728395, - 64'd2947750446693449, 64'd358506668139408, 64'd164866210802549, 64'd10581425453120, - 64'd3100085157486335, 64'd251015876648252, 64'd160926086738718, 64'd13300130662146, - 64'd3198977603974963, 64'd144990905204422, 64'd154784558900806, 64'd15689713641879, - 64'd3245541635063718, 64'd41936768376513, 64'd146639339622086, 64'd17730569029005, - 64'd3241615022546059, - 64'd56758437035189, 64'd136708364113510, 64'd19409222543207},
		'{64'd11799314100150670, 64'd1726645102791665, 64'd334163755354307, 64'd48561971159818, 64'd10952591127214628, 64'd1659711317154405, 64'd323753374549305, 64'd49015407026636, 64'd10139804252581744, 64'd1591020420745462, 64'd312702769499617, 64'd49143758653124, 64'd9361683830509244, 64'd1521154085508429, 64'd301145711237301, 64'd48982853438203, 64'd8618684244533847, 64'd1450635166671628, 64'd289203764829884, 64'd48566108769607, 64'd7911012390371385, 64'd1379931390804498, 64'd276986981713980, 64'd47924616070612, 64'd7238654340870150, 64'd1309458937568988, 64'd264594578586406, 64'd47087228405991, 64'd6601400248267951, 64'd1239585907086178, 64'd252115600567391, 64'd46080650757144, 64'd5998867542649463, 64'd1170635666386360, 64'd239629566695339, 64'd44929532161494, 64'd5430522488407580, 64'd1102890069821280, 64'd227207096129585, 64'd43656558991310, 64'd4895700162747228, 64'd1036592549597817, 64'd214910513727958, 64'd42282548722202, 64'd4393622921895572, 64'd971951073750469, 64'd202794433931221, 64'd40826543611873, 64'd3923417421757894, 64'd909140969912908, 64'd190906322127786, 64'd39305903775323, 64'd3484130260339856, 64'd848307614183701, 64'd179287032890993, 64'd37736399203861, 64'd3074742309396342, 64'd789568985214973, 64'd167971324678882, 64'd36132300332036, 64'd2694181802513566, 64'd733018084392030, 64'd156988350764125, 64'd34506466809278, 64'd2341336246230446, 64'd678725223623238, 64'd146362126320812, 64'd32870434181603, 64'd2015063219899441, 64'd626740182829036, 64'd136111971736398, 64'd31234498233591, 64'd1714200128815726, 64'd577094239712797, 64'd126252932342361, 64'd29607796781994, 64'd1437572973743111, 64'd529802074820183, 64'd116796174867260, 64'd27998388750033},
		'{- 64'd11799314100150724, - 64'd1726645102791664, - 64'd334163755354309, - 64'd48561971159818, - 64'd10952591127214666, - 64'd1659711317154402, - 64'd323753374549306, - 64'd49015407026636, - 64'd10139804252581770, - 64'd1591020420745457, - 64'd312702769499617, - 64'd49143758653124, - 64'd9361683830509258, - 64'd1521154085508422, - 64'd301145711237302, - 64'd48982853438203, - 64'd8618684244533850, - 64'd1450635166671619, - 64'd289203764829885, - 64'd48566108769607, - 64'd7911012390371378, - 64'd1379931390804488, - 64'd276986981713981, - 64'd47924616070612, - 64'd7238654340870134, - 64'd1309458937568976, - 64'd264594578586406, - 64'd47087228405991, - 64'd6601400248267928, - 64'd1239585907086164, - 64'd252115600567391, - 64'd46080650757144, - 64'd5998867542649432, - 64'd1170635666386346, - 64'd239629566695339, - 64'd44929532161494, - 64'd5430522488407544, - 64'd1102890069821265, - 64'd227207096129585, - 64'd43656558991310, - 64'd4895700162747188, - 64'd1036592549597802, - 64'd214910513727958, - 64'd42282548722202, - 64'd4393622921895528, - 64'd971951073750454, - 64'd202794433931221, - 64'd40826543611872, - 64'd3923417421757846, - 64'd909140969912892, - 64'd190906322127786, - 64'd39305903775323, - 64'd3484130260339806, - 64'd848307614183685, - 64'd179287032890993, - 64'd37736399203861, - 64'd3074742309396289, - 64'd789568985214957, - 64'd167971324678882, - 64'd36132300332036, - 64'd2694181802513512, - 64'd733018084392014, - 64'd156988350764125, - 64'd34506466809278, - 64'd2341336246230391, - 64'd678725223623223, - 64'd146362126320812, - 64'd32870434181603, - 64'd2015063219899384, - 64'd626740182829020, - 64'd136111971736398, - 64'd31234498233591, - 64'd1714200128815670, - 64'd577094239712781, - 64'd126252932342361, - 64'd29607796781994, - 64'd1437572973743055, - 64'd529802074820168, - 64'd116796174867260, - 64'd27998388750033}};

	localparam logic signed[63:0] hf[0:1599] = {64'd11750322733056, - 64'd74886045696, - 64'd97475510272, 64'd1163145600, 64'd11675535147008, - 64'd223675695104, - 64'd94927912960, 64'd3450310400, 64'd11527000162304, - 64'd369577066496, - 64'd89903644672, 64'd5625255424, 64'd11306625138688, - 64'd510757699584, - 64'd82525061120, 64'd7624293376, 64'd11017209774080, - 64'd645478023168, - 64'd72958746624, 64'd9393492992, 64'd10662394724352, - 64'd772119461888, - 64'd61409513472, 64'd10888738816, 64'd10246593445888, - 64'd889208700928, - 64'd48114200576, 64'd12075640832, 64'd9774915649536, - 64'd995438755840, - 64'd33335392256, 64'd12929331200, 64'd9253082365952, - 64'd1089685422080, - 64'd17355098112, 64'd13434120192, 64'd8687323185152, - 64'd1171020578816, - 64'd468549088, 64'd13583058944, 64'd8084283981824, - 64'd1238720839680, 64'd17021834240, 64'd13377393664, 64'd7450919436288, - 64'd1292273057792, 64'd34812235776, 64'd12825938944, 64'd6794387128320, - 64'd1331375636480, 64'd52602888192, 64'd11944381440, 64'd6121943728128, - 64'd1355936825344, 64'd70103154688, 64'd10754521088, 64'd5440839614464, - 64'd1366068690944, 64'd87036157952, 64'd9283473408, 64'd4758220308480, - 64'd1362079252480, 64'd103142899712, 64'd7562837504, 64'd4081030266880, - 64'd1344461209600, 64'd118185910272, 64'd5627850240, 64'd3415924277248, - 64'd1313877655552, 64'd131952304128, 64'd3516536576, 64'd2769186455552, - 64'd1271147397120, 64'd144256286720, 64'd1268868992, 64'd2146656190464, - 64'd1217226473472, 64'd154941095936, - 64'd1074052864, 64'd1553664311296, - 64'd1153189150720, 64'd163880353792, - 64'd3470788608, 64'd994978955264, - 64'd1080208654336, 64'd170978902016, - 64'd5880304128, 64'd474761494528, - 64'd999535869952, 64'd176173039616, - 64'd8262667776, - 64'd3467157760, - 64'd912478306304, 64'd179430260736, - 64'd10579685376, - 64'd436849737728, - 64'd820379385856, 64'd180748550144, - 64'd12795478016, - 64'd823205232640, - 64'd724597342208, 64'd180155154432, - 64'd14876981248, - 64'd1161031319552, - 64'd626485559296, 64'd177704992768, - 64'd16794379264, - 64'd1449496936448, - 64'd527373205504, 64'd173478739968, - 64'd18521458688, - 64'd1688426119168, - 64'd428547145728, 64'd167580467200, - 64'd20035887104, - 64'd1878271852544, - 64'd331235688448, 64'd160135168000, - 64'd21319415808, - 64'd2020083630080, - 64'd236593250304, 64'd151286005760, - 64'd22357999616, - 64'd2115466821632, - 64'd145687265280, 64'd141191397376, - 64'd23141857280, - 64'd2166536404992, - 64'd59486650368, 64'd130021974016, - 64'd23665444864, - 64'd2175865061376, 64'd21147623424, 64'd117957582848, - 64'd23927373824, - 64'd2146427207680, 64'd95470043136, 64'd105184174080, - 64'd23930263552, - 64'd2081540276224, 64'd162856026112, 64'd91890761728, - 64'd23680530432, - 64'd1984802586624, 64'd222805360640, 64'd78266564608, - 64'd23188148224, - 64'd1860031348736, 64'd274943770624, 64'd64498094080, - 64'd22466334720, - 64'd1711199354880, 64'd319022366720, 64'd50766598144, - 64'd21531222016, - 64'd1542372982784, 64'd354915614720, 64'd37245579264, - 64'd20401498112, - 64'd1357651378176, 64'd382617223168, 64'd24098566144, - 64'd19098007552, - 64'd1161107603456, 64'd402234900480, 64'd11477163008, - 64'd17643358208, - 64'd956734504960, 64'd413983211520, - 64'd480663840, - 64'd16061496320, - 64'd748392087552, 64'd418175746048, - 64'd11652013056, - 64'd14377304064, - 64'd539760820224, 64'd415215681536, - 64'd21930182656, - 64'd12616183808, - 64'd334299267072, 64'd405585920000, - 64'd31225513984, - 64'd10803657728, - 64'd135206821888, 64'd389838274560, - 64'd39465943040, - 64'd8964982784, 64'd54607884288, 64'd368582164480, - 64'd46597279744, - 64'd7124793856, 64'd232552988672, 64'd342473211904, - 64'd52583174144, - 64'd5306759680, 64'd396373491712, 64'd312201445376, - 64'd57404878848, - 64'd3533280768, 64'd544165625856, 64'd278479634432, - 64'd61060698112, - 64'd1825212288, 64'd674385297408, 64'd242032066560, - 64'd63565250560, - 64'd201625520, 64'd785851154432, 64'd203583389696, - 64'd64948531200, 64'd1320393728, 64'd877741932544, 64'd163848126464, - 64'd65254752256, 64'd2725907968, 64'd949589114880, 64'd123520827392, - 64'd64541057024, 64'd4002252032, 64'd1001264578560, 64'd83267051520, - 64'd62876114944, 64'd5139117568, 64'd1032963883008, 64'd43715047424, - 64'd60338556928, 64'd6128597504, 64'd1045185953792, 64'd5448553984, - 64'd57015418880, 64'd6965194752, 64'd1038709030912, - 64'd30999502848, - 64'd53000454144, 64'd7645795328, 64'd1014563930112, - 64'd65152225280, - 64'd48392486912, 64'd8169603584, 64'd974005207040, - 64'd96592879616, - 64'd43293720576, 64'd8538050048, 64'd918479896576, - 64'd124967968768, - 64'd37808123904, 64'd8754670592, 64'd849595596800, - 64'd149989212160, - 64'd32039831552, 64'd8824955904, 64'd769087504384, - 64'd171434475520, - 64'd26091620352, 64'd8756187136, 64'd678785384448, - 64'd189147660288, - 64'd20063502336, 64'd8557241856, 64'd580580605952, - 64'd203037655040, - 64'd14051398656, 64'd8238396416, 64'd476394389504, - 64'd213076410368, - 64'd8145952256, 64'd7811109888, 64'd368146677760, - 64'd219296038912, - 64'd2431468800, 64'd7287802368, 64'd257726988288, - 64'd221785423872, 64'd3014998784, 64'd6681631744, 64'd146967183360, - 64'd220685877248, 64'd8124414464, 64'd6006267904, 64'd37616291840, - 64'd216186388480, 64'd12836367360, 64'd5275669504, - 64'd68682022912, - 64'd208518463488, 64'd17099527168, 64'd4503869440, - 64'd170409279488, - 64'd197950423040, 64'd20871942144, 64'd3704766720, - 64'd266189127680, - 64'd184781537280, 64'd24121186304, 64'd2891932928, - 64'd354801385472, - 64'd169335980032, 64'd26824353792, 64'd2078429952, - 64'd435192856576, - 64'd151956783104, 64'd28967927808, 64'd1276646016, - 64'd506485309440, - 64'd132999585792, 64'd30547496960, 64'd498147840, - 64'd567980261376, - 64'd112826810368, 64'd31567370240, - 64'd246446752, - 64'd619160862720, - 64'd91801772032, 64'd32040075264, - 64'd947577280, - 64'd659691012096, - 64'd70283206656, 64'd31985752064, - 64'd1596827648, - 64'd689411850240, - 64'd48620093440, 64'd31431479296, - 64'd2186992128, - 64'd708335304704, - 64'd27146878976, 64'd30410520576, - 64'd2712121600, - 64'd716636225536, - 64'd6179153408, 64'd28961515520, - 64'd3167546368, - 64'd714641571840, 64'd13990170624, 64'd27127644160, - 64'd3549882880, - 64'd702818549760, 64'd33094158336, 64'd24955744256, - 64'd3857017344, - 64'd681760456704, 64'd50894602240, 64'd22495436800, - 64'd4088074240, - 64'd652172394496, 64'd67184209920, 64'd19798247424, - 64'd4243367424, - 64'd614854754304, 64'd81788223488, 64'd16916731904, - 64'd4324334080, - 64'd570687094784, 64'd94565449728, 64'd13903649792, - 64'd4333459968, - 64'd520610938880, 64'd105408782336, 64'd10811156480, - 64'd4274186240, - 64'd465612931072, 64'd114245165056, 64'd7690058240, - 64'd4150814208, - 64'd406707765248, 64'd121035022336, 64'd4589113344, - 64'd3968395008, - 64'd344921800704, 64'd125771284480, 64'd1554405120, - 64'd3732619776, - 64'd281277071360, 64'd128477880320, - 64'd1371218304, - 64'd3449700096, - 64'd216776228864, 64'd129207951360, - 64'd4148626176, - 64'd3126251776, - 64'd152388599808, 64'd128041590784, - 64'd6742810112, - 64'd2769174016, - 64'd89037135872, 64'd125083426816, - 64'd9123207168, - 64'd2385533440, - 64'd27586971648, 64'd120459829248, - 64'd11263939584, - 64'd1982449920, 64'd31164805120, 64'd114316001280, - 64'd13143974912, - 64'd1566986880, 64'd86497771520, 64'd106812932096, - 64'd14747205632, - 64'd1146049152, 64'd137775284224, 64'd98124210176, - 64'd16062450688, - 64'd726286848, 64'd184449974272, 64'd88432828416, - 64'd17083383808, - 64'd314008608, 64'd226067693568, 64'd77928062976, - 64'd17808392192, 64'd84895976, 64'd262269779968, 64'd66802278400, - 64'd18240374784, 64'd465024256, 64'd292793942016, 64'd55247974400, - 64'd18386477056, 64'd821517440, 64'd317473587200, 64'd43454877696, - 64'd18257784832, 64'd1150106752, 64'd336235626496, 64'd31607265280, - 64'd17868959744, 64'd1447148672, 64'd349097361408, 64'd19881496576, - 64'd17237856256, 64'd1709648896, 64'd356161716224, 64'd8443739136, - 64'd16385100800, 64'd1935275520, 64'd357611765760, - 64'd2551986688, - 64'd15333640192, 64'd2122361984, 64'd353704181760, - 64'd12965530624, - 64'd14108300288, 64'd2269899264, 64'd344761925632, - 64'd22672025600, - 64'd12735316992, 64'd2377520128, 64'd331166384128, - 64'd31563016192, - 64'd11241880576, 64'd2445471744, 64'd313348784128, - 64'd39547273216, - 64'd9655682048, 64'd2474584064, 64'd291781672960, - 64'd46551339008, - 64'd8004477952, 64'd2466228480, 64'd266969694208, - 64'd52519747584, - 64'd6315674624, 64'd2422271232, 64'd239440838656, - 64'd57415000064, - 64'd4615933440, 64'd2345021440, 64'd209737318400, - 64'd61217263616, - 64'd2930811136, 64'd2237175552, 64'd178407014400, - 64'd63923793920, - 64'd1284432768, 64'd2101758592, 64'd145995038720, - 64'd65548181504, 64'd300799328, 64'd1942062592, 64'd113035845632, - 64'd66119352320, 64'd1804456704, 64'd1761585408, 64'd80045785088, - 64'd65680412672, 64'd3208293632, 64'd1563967872, 64'd47516426240, - 64'd64287309824, 64'd4496413696, 64'd1352933248, 64'd15908431872, - 64'd62007406592, 64'd5655393792, 64'd1132227328, - 64'd14353744896, - 64'd58917916672, 64'd6674364928, 64'd905561792, - 64'd42886389760, - 64'd55104299008, 64'd7545052160, 64'd676560192, - 64'd69350219776, - 64'd50658578432, 64'd8261770752, 64'd448708736, - 64'd93453279232, - 64'd45677682688, 64'd8821388288, 64'd225310528, - 64'd114952921088, - 64'd40261754880, 64'd9223249920, 64'd9445386, - 64'd133657059328, - 64'd34512523264, 64'd9469064192, - 64'd196065376, - 64'd149424504832, - 64'd28531697664, 64'd9562771456, - 64'd388688512, - 64'd162164637696, - 64'd22419496960, 64'd9510370304, - 64'd566202624, - 64'd171836260352, - 64'd16273199104, 64'd9319736320, - 64'd726716288, - 64'd178445762560, - 64'd10185863168, 64'd9000410112, - 64'd868680512, - 64'd182044835840, - 64'd4245144320, 64'd8563378688, - 64'd990894976, - 64'd182727376896, 64'd1467744128, 64'd8020840960, - 64'd1092509440, - 64'd180626096128, 64'd6878921728, 64'd7385970688, - 64'd1173019392, - 64'd175908651008, 64'd11922582528, 64'd6672670208, - 64'd1232257024, - 64'd168773468160, 64'd16541582336, 64'd5895333376, - 64'd1270377728, - 64'd159445270528, 64'd20687863808, 64'd5068605952, - 64'd1287841920, - 64'd148170473472, 64'd24322734080, 64'd4207155456, - 64'd1285393664, - 64'd135212507136, 64'd27416981504, 64'd3325454848, - 64'd1264035968, - 64'd120846983168, 64'd29950849024, 64'd2437575680, - 64'd1225004032, - 64'd105357090816, 64'd31913873408, 64'd1556998656, - 64'd1169734528, - 64'd89028984832, 64'd33304588288, 64'd696442752, - 64'd1099835648, - 64'd72147369984, 64'd34130106368, - 64'd132287264, - 64'd1017054656, - 64'd54991368192, 64'd34405605376, - 64'd918431360, - 64'd923245120, - 64'd37830623232, 64'd34153697280, - 64'd1652383616, - 64'd820334336, - 64'd20921751552, 64'd33403754496, - 64'd2325779200, - 64'd710291456, - 64'd4505156096, 64'd32191121408, - 64'd2931558144, - 64'd595095744, 64'd11197762560, 64'd30556315648, - 64'd3464007424, - 64'd476707168, 64'd25986973696, 64'd28544169984, - 64'd3918779648, - 64'd357038080, 64'd39685758976, 64'd26202953728, - 64'd4292892928, - 64'd237927136, 64'd52142219264, 64'd23583496192, - 64'd4584708096, - 64'd121115528, 64'd63230308352, 64'd20738297856, - 64'd4793888256, - 64'd8225954, 64'd72850481152, 64'd17720678400, - 64'd4921340416, 64'd99255800, 64'd80929882112, 64'd14583931904, - 64'd4969142784, 64'd199996272, 64'd87422132224, 64'd11380551680, - 64'd4940455936, 64'd292826784, 64'd92306718720, 64'd8161475072, - 64'd4839424000, 64'd376752768, 64'd95588089856, 64'd4975407104, - 64'd4671066112, 64'd450960128, 64'd97294360576, 64'd1868203392, - 64'd4441157632, 64'd514818656, 64'd97475715072, - 64'd1117672704, - 64'd4156110592, 64'd567882368, 64'd96202661888, - 64'd3943618816, - 64'd3822844416, 64'd609887296, 64'd93563920384, - 64'd6575279616, - 64'd3448660480, 64'd640746624, 64'd89664290816, - 64'd8982853632, - 64'd3041114624, 64'd660543296, 64'd84622270464, - 64'd11141313536, - 64'd2607892992, 64'd669520576, 64'd78567653376, - 64'd13030548480, - 64'd2156690432, 64'd668070912, 64'd71639048192, - 64'd14635427840, - 64'd1695096320, 64'd656722496, 64'd63981359104, - 64'd15945781248, - 64'd1230487168, 64'd636125120, 64'd55743389696, - 64'd16956310528, - 64'd769926784, 64'd607034560, 64'd47075373056, - 64'd17666437120, - 64'd320076672, 64'd570296128, 64'd38126714880, - 64'd18080073728, 64'd112883712, 64'd526827904, 64'd29043789824, - 64'd18205360128, 64'd523325280, 64'd477603552, 64'd19967913984, - 64'd18054326272, 64'd906226560, 64'd423635072, 64'd11033488384, - 64'd17642536960, 64'd1257218688, 64'd365956000, 64'd2366337280, - 64'd16988678144, 64'd1572619008, 64'd305604928, - 64'd5917753856, - 64'd16114135040, 64'd1849452416, 64'd243609840, - 64'd13714274304, - 64'd15042542592, 64'd2085461632, 64'd180973392, - 64'd20930994176, - 64'd13799323648, 64'd2279105536, 64'd118659216, - 64'd27488749568, - 64'd12411227136, 64'd2429548288, 64'd57579436, - 64'd33321981952, - 64'd10905863168, 64'd2536636160, - 64'd1416332, - 64'd38379057152, - 64'd9311252480, 64'd2600868864, - 64'd57550620, - 64'd42622369792, - 64'd7655389184, 64'd2623358208, - 64'd110126160, - 64'd46028210176, - 64'd5965828096, 64'd2605783808, - 64'd158532384, - 64'd48586457088, - 64'd4269294080, 64'd2550340352, - 64'd202250272, - 64'd50300067840, - 64'd2591324928, 64'd2459678464, - 64'd240855680, - 64'd51184402432, - 64'd955949696, 64'd2336845568, - 64'd274021024, - 64'd51266400256, 64'd614595456, 64'd2185219584, - 64'd301515488, - 64'd50583621632, 64'd2100111616, 64'd2008443648, - 64'd323203744, - 64'd49183158272, 64'd3482639104, 64'd1810359040, - 64'd339043456, - 64'd47120510976, 64'd4746615808, 64'd1594937984, - 64'd349081184, - 64'd44458311680, 64'd5878992384, 64'd1366218752, - 64'd353447680, - 64'd41265094656, 64'd6869306880, 64'd1128242432, - 64'd352351648, - 64'd37613957120, 64'd7709711872, 64'd884992128, - 64'd346072928, - 64'd33581264896, 64'd8394967040, 64'd640337408, - 64'd334954976, - 64'd29245374464, 64'd8922391552, 64'd397981504, - 64'd319396544, - 64'd24685348864, 64'd9291779072, 64'd161414864, - 64'd299843200, - 64'd19979759616, 64'd9505280000, - 64'd66126916, - 64'd276778400, - 64'd15205549056, 64'd9567258624, - 64'd281698560, - 64'd250714416, - 64'd10436952064, 64'd9484120064, - 64'd482674976, - 64'd222183376, - 64'd5744536576, 64'd9264114688, - 64'd666774848, - 64'd191728400, - 64'd1194323712, 64'd8917130240, - 64'd832077888, - 64'd159894976, 64'd3152969728, 64'd8454461440, - 64'd977035904, - 64'd127222720, 64'd7242577408, 64'd7888576000, - 64'd1100477824, - 64'd94237664, 64'd11026210816, 64'd7232873984, - 64'd1201609088, - 64'd61445076, 64'd14462461952, 64'd6501441024, - 64'd1280004864, - 64'd29322966, 64'd17517086720, 64'd5708808704, - 64'd1335598848, 64'd1683714, 64'd20163170304, 64'd4869714432, - 64'd1368667008, 64'd31168090, 64'd22381168640, 64'd3998873344, - 64'd1379806336, 64'd58765564, 64'd24158840832, 64'd3110761984, - 64'd1369911040, 64'd84157200, 64'd25491087360, 64'd2219412736, - 64'd1340144896, 64'd107072248, 64'd26379669504, 64'd1338227968, - 64'd1291910528, 64'd127289848, 64'd26832861184, 64'd479810912, - 64'd1226817152, 64'd144639904, 64'd26865000448, - 64'd344182848, - 64'd1146647168, 64'd159003152, 64'd26495991808, - 64'd1123172992, - 64'd1053320256, 64'd170310480, 64'd25750740992, - 64'd1847759488, - 64'd948859328, 64'd178541536, 64'd24658536448, - 64'd2509805568, - 64'd835354880, 64'd183722656, 64'd23252410368, - 64'd3102496768, - 64'd714930688, 64'd185924240, 64'd21568458752, - 64'd3620379904, - 64'd589710656, 64'd185257568, 64'd19645161472, - 64'd4059376128, - 64'd461787456, 64'd181871168, 64'd17522694144, - 64'd4416777216, - 64'd333192640, 64'd175946800, 64'd15242254336, - 64'd4691217920, - 64'd205869584, 64'd167695168, 64'd12845386752, - 64'd4882632192, - 64'd81648800, 64'd157351376, 64'd10373361664, - 64'd4992191488, 64'd37773780, 64'd145170240, 64'd7866569728, - 64'd5022226432, 64'd150855536, 64'd131421576, 64'd5363962880, - 64'd4976137216, 64'd256222624, 64'd116385472, 64'd2902548480, - 64'd4858291712, 64'd352682304, 64'd100347592, 64'd516930752, - 64'd4673911808, 64'd439231904, 64'd83594680, - 64'd1761086592, - 64'd4428957184, 64'd515064448, 64'd66410244, - 64'd3902837248, - 64'd4129998080, 64'd579571264, 64'd49070508, - 64'd5883067392, - 64'd3784090880, 64'd632341440, 64'd31840648, - 64'd7680145408, - 64'd3398648064, 64'd673158400, 64'd14971387, - 64'd9276208128, - 64'd2981311488, 64'd701993600, - 64'd1304030, - 64'd10657245184, - 64'd2539827456, 64'd718998080, - 64'd16772460, - 64'd11813120000, - 64'd2081926272, 64'd724491200, - 64'd31243058, - 64'd12737531904, - 64'd1615208960, 64'd718948160, - 64'd44549036, - 64'd13427928064, - 64'd1147039616, 64'd702985152, - 64'd56548972, - 64'd13885356032, - 64'd684448128, 64'd677343360, - 64'd67127696, - 64'd14114276352, - 64'd234041408, 64'd642872064, - 64'd76196728, - 64'd14122331136, 64'd198074304, 64'd600510656, - 64'd83694304, - 64'd13920076800, 64'd606359808, 64'd551270464, - 64'd89584992, - 64'd13520683008, 64'd985897920, 64'd496216000, - 64'd93858968, - 64'd12939616256, 64'd1332436736, 64'd436446816, - 64'd96530904, - 64'd12194294784, 64'd1642420224, 64'd373079424, - 64'd97638568, - 64'd11303736320, 64'd1913007616, 64'd307229664, - 64'd97241152, - 64'd10288197632, 64'd2142081536, 64'd239996480, - 64'd95417360, - 64'd9168815104, 64'd2328243456, 64'd172446144, - 64'd92263288, - 64'd7967245824, 64'd2470800640, 64'd105598096, - 64'd87890152, - 64'd6705322496, 64'd2569741824, 64'd40412068, - 64'd82421920, - 64'd5404718592, 64'd2625704960, - 64'd22223332, - 64'd75992832, - 64'd4086636288, 64'd2639935744, - 64'd81500376, - 64'd68744912, - 64'd2771511296, 64'd2614240000, - 64'd136700320, - 64'd60825504, - 64'd1478748032, 64'd2550929664, - 64'd187199744, - 64'd52384792, - 64'd226480688, 64'd2452763904, - 64'd232475280, - 64'd43573456, 64'd968635264, 64'd2322886656, - 64'd272106496, - 64'd34540396, 64'd2091598976, 64'd2164761856, - 64'd305777152, - 64'd25430600, 64'd3129207040, 64'd1982104576, - 64'd333274944, - 64'd16383198, 64'd4070163456, 64'd1778816128, - 64'd354489568, - 64'd7529658, 64'd4905154048, 64'd1558915200, - 64'd369409440, 64'd1007791, 64'd5626890240, 64'd1326473344, - 64'd378117120, 64'd9117525, 64'd6230119424, 64'd1085551744, - 64'd380783488, 64'd16699677, 64'd6711604224, 64'd840141184, - 64'd377660960, 64'd23667050, 64'd7070073344, 64'd594106176, - 64'd369075840, 64'd29945802, 64'd7306144768, 64'd351133920, - 64'd355419776, 64'd35475892, 64'd7422226432, 64'd114687632, - 64'd337140928, 64'd40211324, 64'd7422393344, - 64'd112033768, - 64'd314734464, 64'd44120116, 64'd7312246272, - 64'd326130592, - 64'd288732960, 64'd47184140, 64'd7098754048, - 64'd525031008, - 64'd259696704, 64'd49398688, 64'd6790086144, - 64'd706513344, - 64'd228203968, 64'd50771912, 64'd6395430400, - 64'd868722176, - 64'd194841632, 64'd51324076, 64'd5924809216, - 64'd1010178368, - 64'd160195936, 64'd51086660, 64'd5388889600, - 64'd1129782656, - 64'd124843896, 64'd50101372, 64'd4798793216, - 64'd1226813696, - 64'd89345112, 64'd48419008, 64'd4165909504, - 64'd1300920576, - 64'd54234316, 64'd46098272, 64'd3501712896, - 64'd1352110080, - 64'd20014620, 64'd43204520, 64'd2817588480, - 64'd1380729216, 64'd12848429, 64'd39808472, 64'd2124667904, - 64'd1387443840, 64'd43931956, 64'd35984880, 64'd1433674624, - 64'd1373212928, 64'd72859984, 64'd31811254, 64'd754785408, - 64'd1339260800, 64'd99306744, 64'd27366544, 64'd97505080, - 64'd1287045248, 64'd122999096, 64'd22729924, - 64'd529442272, - 64'd1218225408, 64'd143718064, 64'd17979584, - 64'd1118205056, - 64'd1134626816, 64'd161299408, 64'd13191634, - 64'd1661879040, - 64'd1038206528, 64'd175633520, 64'd8439054, - 64'd2154563328, - 64'd931017408, 64'd186664304, 64'd3790776, - 64'd2591400960, - 64'd815173248, 64'd194387520, - 64'd689153, - 64'd2968599296, - 64'd692814272, 64'd198848272, - 64'd4942285, - 64'd3283435520, - 64'd566074048, 64'd200137952, - 64'd8916367, - 64'd3534245632, - 64'd437048064, 64'd198390720, - 64'd12565821, - 64'd3720397056, - 64'd307764608, 64'd193779344, - 64'd15852098, - 64'd3842249728, - 64'd180157664, 64'd186510832, - 64'd18743908, - 64'd3901101056, - 64'd56042756, 64'd176821664, - 64'd21217340, - 64'd3899122432, 64'd62904204, 64'd164972880, - 64'd23255856, - 64'd3839284480, 64'd175165168, 64'd151244992, - 64'd24850182, - 64'd3725274112, 64'd279394848, 64'd135932864, - 64'd25998096, - 64'd3561405184, 64'd374432320, 64'd119340704, - 64'd26704114, - 64'd3352523520, 64'd459309536, 64'd101776976, - 64'd26979106, - 64'd3103910400, 64'd533256096, 64'd83549712, - 64'd26839824, - 64'd2821182208, 64'd595701440, 64'd64961900, - 64'd26308364, - 64'd2510190592, 64'd646273472, 64'd46307240, - 64'd25411584, - 64'd2176924160, 64'd684794560, 64'd27866232, - 64'd24180474, - 64'd1827413632, 64'd711274816, 64'd9902631, - 64'd22649494, - 64'd1467639296, 64'd725902784, - 64'd7339646, - 64'd20855898, - 64'd1103444736, 64'd729034112, - 64'd23639200, - 64'd18839040, - 64'd740456960, 64'd721178112, - 64'd38799348, - 64'd16639687, - 64'd384012864, 64'd702982656, - 64'd52649852, - 64'd14299354, - 64'd39094080, 64'd675218176, - 64'd65048160, - 64'd11859640, 64'd289729920, 64'd638759936, - 64'd75880208, - 64'd9361610, 64'd598349824, 64'd594570112, - 64'd85060728, - 64'd6845214, 64'd883155264, 64'd543679424, - 64'd92533104, - 64'd4348738, 64'd1141064448, 64'd487168128, - 64'd98268856, - 64'd1908327, 64'd1369544192, 64'd426148000, - 64'd102266704, 64'd442460, 64'd1566621312, 64'd361743968, - 64'd104551240, 64'd2673014, 64'd1730884992, 64'd295076864, - 64'd105171344, 64'd4755996, 64'd1861479936, 64'd227247040, - 64'd104198272, 64'd6667580, 64'd1958092800, 64'd159318864, - 64'd101723504, 64'd8387642, 64'd2020930560, 64'd92306752, - 64'd97856440, 64'd9899874, 64'd2050692096, 64'd27162426, - 64'd92721856, 64'd11191850, 64'd2048534272, - 64'd35236140, - 64'd86457360, 64'd12255013, 64'd2016032128, - 64'd94094240, - 64'd79210688, 64'd13084626, 64'd1955136000, - 64'd148708208, - 64'd71137032, 64'd13679647, 64'd1868123776, - 64'd198471504, - 64'd62396380, 64'd14042576, 64'd1757551104, - 64'd242878960, - 64'd53150888, 64'd14179239, 64'd1626200704, - 64'd281529472, - 64'd43562384, 64'd14098545, 64'd1477029504, - 64'd314126912, - 64'd33789972, 64'd13812199, 64'd1313116032, - 64'd340479424, - 64'd23987790, 64'd13334403, 64'd1137609600, - 64'd360497184, - 64'd14302971, 64'd12681513, 64'd953679040, - 64'd374188960, - 64'd4873792, 64'd11871698, 64'd764465536, - 64'd381657056, 64'd4171960, 64'd10924582, 64'd573036992, - 64'd383091392, 64'd12718370, 64'd9860880, 64'd382345600, - 64'd378762368, 64'd20662552, 64'd8702040, 64'd195190160, - 64'd369012896, 64'd27915546, 64'd7469884, 64'd14181419, - 64'd354250016, 64'd34402964, 64'd6186271, - 64'd158287360, - 64'd334935488, 64'd40065392, 64'd4872768, - 64'd320065568, - 64'd311576480, 64'd44858552, 64'd3550343, - 64'd469265472, - 64'd284715680, 64'd48753232, 64'd2239082, - 64'd604277632, - 64'd254921632, 64'd51734980, 64'd957937, - 64'd723781120, - 64'd222779008, 64'd53803616, - 64'd275508, - 64'd826749504, - 64'd188879088, 64'd54972532, - 64'd1445224, - 64'd912451840, - 64'd153810704, 64'd55267860, - 64'd2536908, - 64'd980448896, - 64'd118151560, 64'd54727440, - 64'd3538106, - 64'd1030586048, - 64'd82460240, 64'd53399712, - 64'd4438312, - 64'd1062981504, - 64'd47268804, 64'd51342476, - 64'd5229027, - 64'd1078011520, - 64'd13076129, 64'd48621572, - 64'd5903792, - 64'd1076292224, 64'd19657844, 64'd45309532, - 64'd6458186, - 64'd1058658880, 64'd50517104, 64'd41484160, - 64'd6889785, - 64'd1026142976, 64'd79133616, 64'd37227136, - 64'd7198112, - 64'd979947392, 64'd105190464, 64'd32622598, - 64'd7384546, - 64'd921419904, 64'd128424112, 64'd27755788, - 64'd7452206, - 64'd852026816, 64'd148625712, 64'd22711724, - 64'd7405830, - 64'd773324672, 64'd165641600, 64'd17573944, - 64'd7251620, - 64'd686933440, 64'd179372880, 64'd12423344, - 64'd6997082, - 64'd594508800, 64'd189774240, 64'd7337101, - 64'd6650849, - 64'd497716160, 64'd196852080, 64'd2387700, - 64'd6222502, - 64'd398205440, 64'd200661888, - 64'd2357908, - 64'd5722375, - 64'd297587040, 64'd201305008, - 64'd6839042, - 64'd5161374, - 64'd197410032, 64'd198924992, - 64'd11001883, - 64'd4550779, - 64'd99142048, 64'd193703360, - 64'd14799945, - 64'd3902064, - 64'd4151368, 64'd185855120, - 64'd18194412, - 64'd3226714, 64'd86308584, 64'd175623888, - 64'd21154344, - 64'd2536054, 64'd171112320, 64'd163276960, - 64'd23656752, - 64'd1841090, 64'd249272832, 64'd149100128, - 64'd25686564, - 64'd1152360, 64'd319949568, 64'd133392576, - 64'd27236456, - 64'd479799, 64'd382453888, 64'd116461768, - 64'd28306596, 64'd167379, 64'd436251808, 64'd98618496, - 64'd28904270, 64'd780780, 64'd480964704, 64'd80172080, - 64'd29043436, 64'd1352921, 64'd516367168, 64'd61425856, - 64'd28744196, 64'd1877293, 64'd542383168, 64'd42672952, - 64'd28032188, 64'd2348411, 64'd559079808, 64'd24192414, - 64'd26937954, 64'd2761848, 64'd566659456, 64'd6245758, - 64'd25496234, 64'd3114246, 64'd565450240, - 64'd10926079, - 64'd23745258, 64'd3403320, 64'd555894976, - 64'd27105328, - 64'd21726004, 64'd3627834, 64'd538539328, - 64'd42099500, - 64'd19481452, 64'd3787572, 64'd514018272, - 64'd55743024, - 64'd17055856, 64'd3883292, 64'd483042688, - 64'd67898416, - 64'd14494022, 64'd3916666, 64'd446385088, - 64'd78456944, - 64'd11840614, 64'd3890212, 64'd404864960, - 64'd87338888, - 64'd9139497, 64'd3807215, 64'd359334560, - 64'd94493272, - 64'd6433125, 64'd3671643, 64'd310664480, - 64'd99897296, - 64'd3761978, 64'd3488053, 64'd259729920, - 64'd103555248, - 64'd1164054, 64'd3261495, 64'd207397392, - 64'd105497184, 64'd1325572, 64'd2997414, 64'd154512336, - 64'd105777200, 64'd3675132, 64'd2701548, 64'd101887520, - 64'd104471472, 64'd5856476, 64'd2379832, 64'd50292516, - 64'd101676088, 64'd7845314, 64'd2038298, 64'd444425, - 64'd97504608, 64'd9621392, 64'd1682980, - 64'd47000308, - 64'd92085560, 64'd11168599, 64'd1319826, - 64'd91452696, - 64'd85559808, 64'd12475003, 64'd954611, - 64'd132396688, - 64'd78077848, 64'd13532828, 64'd592865, - 64'd169393344, - 64'd69797112, 64'd14338368, 64'd239796, - 64'd202083600, - 64'd60879308, 64'd14891849, - 64'd99768, - 64'd230189776, - 64'd51487776, 64'd15197229, - 64'd421433, - 64'd253515744, - 64'd41785008, 64'd15261965, - 64'd721283, - 64'd271945920, - 64'd31930268, 64'd15096727, - 64'd995915, - 64'd285443040, - 64'd22077376, 64'd14715092, - 64'd1242467, - 64'd294044992, - 64'd12372688, 64'd14133192, - 64'd1458633, - 64'd297860608, - 64'd2953286, 64'd13369359, - 64'd1642668, - 64'd297064512, 64'd6054622, 64'd12443741, - 64'd1793389, - 64'd291891584, 64'd14537041, 64'd11377918, - 64'd1910169, - 64'd282630240, 64'd22393300, 64'd10194511, - 64'd1992911, - 64'd269615840, 64'd29536902, 64'd8916792, - 64'd2042032, - 64'd253223232, 64'd35896124, 64'd7568313, - 64'd2058426};

	localparam logic signed[63:0] hb[0:1599] = {64'd11750322733056, 64'd74886045696, - 64'd97475510272, - 64'd1163145600, 64'd11675535147008, 64'd223675695104, - 64'd94927912960, - 64'd3450310400, 64'd11527000162304, 64'd369577066496, - 64'd89903644672, - 64'd5625255424, 64'd11306625138688, 64'd510757699584, - 64'd82525061120, - 64'd7624293376, 64'd11017209774080, 64'd645478023168, - 64'd72958746624, - 64'd9393492992, 64'd10662394724352, 64'd772119461888, - 64'd61409513472, - 64'd10888738816, 64'd10246593445888, 64'd889208700928, - 64'd48114200576, - 64'd12075640832, 64'd9774915649536, 64'd995438755840, - 64'd33335392256, - 64'd12929331200, 64'd9253082365952, 64'd1089685422080, - 64'd17355098112, - 64'd13434120192, 64'd8687323185152, 64'd1171020578816, - 64'd468549088, - 64'd13583058944, 64'd8084283981824, 64'd1238720839680, 64'd17021834240, - 64'd13377393664, 64'd7450919436288, 64'd1292273057792, 64'd34812235776, - 64'd12825938944, 64'd6794387128320, 64'd1331375636480, 64'd52602888192, - 64'd11944381440, 64'd6121943728128, 64'd1355936825344, 64'd70103154688, - 64'd10754521088, 64'd5440839614464, 64'd1366068690944, 64'd87036157952, - 64'd9283473408, 64'd4758220308480, 64'd1362079252480, 64'd103142899712, - 64'd7562837504, 64'd4081030266880, 64'd1344461209600, 64'd118185910272, - 64'd5627850240, 64'd3415924277248, 64'd1313877655552, 64'd131952304128, - 64'd3516536576, 64'd2769186455552, 64'd1271147397120, 64'd144256286720, - 64'd1268868992, 64'd2146656190464, 64'd1217226473472, 64'd154941095936, 64'd1074052864, 64'd1553664311296, 64'd1153189150720, 64'd163880353792, 64'd3470788608, 64'd994978955264, 64'd1080208654336, 64'd170978902016, 64'd5880304128, 64'd474761494528, 64'd999535869952, 64'd176173039616, 64'd8262667776, - 64'd3467157760, 64'd912478306304, 64'd179430260736, 64'd10579685376, - 64'd436849737728, 64'd820379385856, 64'd180748550144, 64'd12795478016, - 64'd823205232640, 64'd724597342208, 64'd180155154432, 64'd14876981248, - 64'd1161031319552, 64'd626485559296, 64'd177704992768, 64'd16794379264, - 64'd1449496936448, 64'd527373205504, 64'd173478739968, 64'd18521458688, - 64'd1688426119168, 64'd428547145728, 64'd167580467200, 64'd20035887104, - 64'd1878271852544, 64'd331235688448, 64'd160135168000, 64'd21319415808, - 64'd2020083630080, 64'd236593250304, 64'd151286005760, 64'd22357999616, - 64'd2115466821632, 64'd145687265280, 64'd141191397376, 64'd23141857280, - 64'd2166536404992, 64'd59486650368, 64'd130021974016, 64'd23665444864, - 64'd2175865061376, - 64'd21147623424, 64'd117957582848, 64'd23927373824, - 64'd2146427207680, - 64'd95470043136, 64'd105184174080, 64'd23930263552, - 64'd2081540276224, - 64'd162856026112, 64'd91890761728, 64'd23680530432, - 64'd1984802586624, - 64'd222805360640, 64'd78266564608, 64'd23188148224, - 64'd1860031348736, - 64'd274943770624, 64'd64498094080, 64'd22466334720, - 64'd1711199354880, - 64'd319022366720, 64'd50766598144, 64'd21531222016, - 64'd1542372982784, - 64'd354915614720, 64'd37245579264, 64'd20401498112, - 64'd1357651378176, - 64'd382617223168, 64'd24098566144, 64'd19098007552, - 64'd1161107603456, - 64'd402234900480, 64'd11477163008, 64'd17643358208, - 64'd956734504960, - 64'd413983211520, - 64'd480663840, 64'd16061496320, - 64'd748392087552, - 64'd418175746048, - 64'd11652013056, 64'd14377304064, - 64'd539760820224, - 64'd415215681536, - 64'd21930182656, 64'd12616183808, - 64'd334299267072, - 64'd405585920000, - 64'd31225513984, 64'd10803657728, - 64'd135206821888, - 64'd389838274560, - 64'd39465943040, 64'd8964982784, 64'd54607884288, - 64'd368582164480, - 64'd46597279744, 64'd7124793856, 64'd232552988672, - 64'd342473211904, - 64'd52583174144, 64'd5306759680, 64'd396373491712, - 64'd312201445376, - 64'd57404878848, 64'd3533280768, 64'd544165625856, - 64'd278479634432, - 64'd61060698112, 64'd1825212288, 64'd674385297408, - 64'd242032066560, - 64'd63565250560, 64'd201625520, 64'd785851154432, - 64'd203583389696, - 64'd64948531200, - 64'd1320393728, 64'd877741932544, - 64'd163848126464, - 64'd65254752256, - 64'd2725907968, 64'd949589114880, - 64'd123520827392, - 64'd64541057024, - 64'd4002252032, 64'd1001264578560, - 64'd83267051520, - 64'd62876114944, - 64'd5139117568, 64'd1032963883008, - 64'd43715047424, - 64'd60338556928, - 64'd6128597504, 64'd1045185953792, - 64'd5448553984, - 64'd57015418880, - 64'd6965194752, 64'd1038709030912, 64'd30999502848, - 64'd53000454144, - 64'd7645795328, 64'd1014563930112, 64'd65152225280, - 64'd48392486912, - 64'd8169603584, 64'd974005207040, 64'd96592879616, - 64'd43293720576, - 64'd8538050048, 64'd918479896576, 64'd124967968768, - 64'd37808123904, - 64'd8754670592, 64'd849595596800, 64'd149989212160, - 64'd32039831552, - 64'd8824955904, 64'd769087504384, 64'd171434475520, - 64'd26091620352, - 64'd8756187136, 64'd678785384448, 64'd189147660288, - 64'd20063502336, - 64'd8557241856, 64'd580580605952, 64'd203037655040, - 64'd14051398656, - 64'd8238396416, 64'd476394389504, 64'd213076410368, - 64'd8145952256, - 64'd7811109888, 64'd368146677760, 64'd219296038912, - 64'd2431468800, - 64'd7287802368, 64'd257726988288, 64'd221785423872, 64'd3014998784, - 64'd6681631744, 64'd146967183360, 64'd220685877248, 64'd8124414464, - 64'd6006267904, 64'd37616291840, 64'd216186388480, 64'd12836367360, - 64'd5275669504, - 64'd68682022912, 64'd208518463488, 64'd17099527168, - 64'd4503869440, - 64'd170409279488, 64'd197950423040, 64'd20871942144, - 64'd3704766720, - 64'd266189127680, 64'd184781537280, 64'd24121186304, - 64'd2891932928, - 64'd354801385472, 64'd169335980032, 64'd26824353792, - 64'd2078429952, - 64'd435192856576, 64'd151956783104, 64'd28967927808, - 64'd1276646016, - 64'd506485309440, 64'd132999585792, 64'd30547496960, - 64'd498147840, - 64'd567980261376, 64'd112826810368, 64'd31567370240, 64'd246446752, - 64'd619160862720, 64'd91801772032, 64'd32040075264, 64'd947577280, - 64'd659691012096, 64'd70283206656, 64'd31985752064, 64'd1596827648, - 64'd689411850240, 64'd48620093440, 64'd31431479296, 64'd2186992128, - 64'd708335304704, 64'd27146878976, 64'd30410520576, 64'd2712121600, - 64'd716636225536, 64'd6179153408, 64'd28961515520, 64'd3167546368, - 64'd714641571840, - 64'd13990170624, 64'd27127644160, 64'd3549882880, - 64'd702818549760, - 64'd33094158336, 64'd24955744256, 64'd3857017344, - 64'd681760456704, - 64'd50894602240, 64'd22495436800, 64'd4088074240, - 64'd652172394496, - 64'd67184209920, 64'd19798247424, 64'd4243367424, - 64'd614854754304, - 64'd81788223488, 64'd16916731904, 64'd4324334080, - 64'd570687094784, - 64'd94565449728, 64'd13903649792, 64'd4333459968, - 64'd520610938880, - 64'd105408782336, 64'd10811156480, 64'd4274186240, - 64'd465612931072, - 64'd114245165056, 64'd7690058240, 64'd4150814208, - 64'd406707765248, - 64'd121035022336, 64'd4589113344, 64'd3968395008, - 64'd344921800704, - 64'd125771284480, 64'd1554405120, 64'd3732619776, - 64'd281277071360, - 64'd128477880320, - 64'd1371218304, 64'd3449700096, - 64'd216776228864, - 64'd129207951360, - 64'd4148626176, 64'd3126251776, - 64'd152388599808, - 64'd128041590784, - 64'd6742810112, 64'd2769174016, - 64'd89037135872, - 64'd125083426816, - 64'd9123207168, 64'd2385533440, - 64'd27586971648, - 64'd120459829248, - 64'd11263939584, 64'd1982449920, 64'd31164805120, - 64'd114316001280, - 64'd13143974912, 64'd1566986880, 64'd86497771520, - 64'd106812932096, - 64'd14747205632, 64'd1146049152, 64'd137775284224, - 64'd98124210176, - 64'd16062450688, 64'd726286848, 64'd184449974272, - 64'd88432828416, - 64'd17083383808, 64'd314008608, 64'd226067693568, - 64'd77928062976, - 64'd17808392192, - 64'd84895976, 64'd262269779968, - 64'd66802278400, - 64'd18240374784, - 64'd465024256, 64'd292793942016, - 64'd55247974400, - 64'd18386477056, - 64'd821517440, 64'd317473587200, - 64'd43454877696, - 64'd18257784832, - 64'd1150106752, 64'd336235626496, - 64'd31607265280, - 64'd17868959744, - 64'd1447148672, 64'd349097361408, - 64'd19881496576, - 64'd17237856256, - 64'd1709648896, 64'd356161716224, - 64'd8443739136, - 64'd16385100800, - 64'd1935275520, 64'd357611765760, 64'd2551986688, - 64'd15333640192, - 64'd2122361984, 64'd353704181760, 64'd12965530624, - 64'd14108300288, - 64'd2269899264, 64'd344761925632, 64'd22672025600, - 64'd12735316992, - 64'd2377520128, 64'd331166384128, 64'd31563016192, - 64'd11241880576, - 64'd2445471744, 64'd313348784128, 64'd39547273216, - 64'd9655682048, - 64'd2474584064, 64'd291781672960, 64'd46551339008, - 64'd8004477952, - 64'd2466228480, 64'd266969694208, 64'd52519747584, - 64'd6315674624, - 64'd2422271232, 64'd239440838656, 64'd57415000064, - 64'd4615933440, - 64'd2345021440, 64'd209737318400, 64'd61217263616, - 64'd2930811136, - 64'd2237175552, 64'd178407014400, 64'd63923793920, - 64'd1284432768, - 64'd2101758592, 64'd145995038720, 64'd65548181504, 64'd300799328, - 64'd1942062592, 64'd113035845632, 64'd66119352320, 64'd1804456704, - 64'd1761585408, 64'd80045785088, 64'd65680412672, 64'd3208293632, - 64'd1563967872, 64'd47516426240, 64'd64287309824, 64'd4496413696, - 64'd1352933248, 64'd15908431872, 64'd62007406592, 64'd5655393792, - 64'd1132227328, - 64'd14353744896, 64'd58917916672, 64'd6674364928, - 64'd905561792, - 64'd42886389760, 64'd55104299008, 64'd7545052160, - 64'd676560192, - 64'd69350219776, 64'd50658578432, 64'd8261770752, - 64'd448708736, - 64'd93453279232, 64'd45677682688, 64'd8821388288, - 64'd225310528, - 64'd114952921088, 64'd40261754880, 64'd9223249920, - 64'd9445386, - 64'd133657059328, 64'd34512523264, 64'd9469064192, 64'd196065376, - 64'd149424504832, 64'd28531697664, 64'd9562771456, 64'd388688512, - 64'd162164637696, 64'd22419496960, 64'd9510370304, 64'd566202624, - 64'd171836260352, 64'd16273199104, 64'd9319736320, 64'd726716288, - 64'd178445762560, 64'd10185863168, 64'd9000410112, 64'd868680512, - 64'd182044835840, 64'd4245144320, 64'd8563378688, 64'd990894976, - 64'd182727376896, - 64'd1467744128, 64'd8020840960, 64'd1092509440, - 64'd180626096128, - 64'd6878921728, 64'd7385970688, 64'd1173019392, - 64'd175908651008, - 64'd11922582528, 64'd6672670208, 64'd1232257024, - 64'd168773468160, - 64'd16541582336, 64'd5895333376, 64'd1270377728, - 64'd159445270528, - 64'd20687863808, 64'd5068605952, 64'd1287841920, - 64'd148170473472, - 64'd24322734080, 64'd4207155456, 64'd1285393664, - 64'd135212507136, - 64'd27416981504, 64'd3325454848, 64'd1264035968, - 64'd120846983168, - 64'd29950849024, 64'd2437575680, 64'd1225004032, - 64'd105357090816, - 64'd31913873408, 64'd1556998656, 64'd1169734528, - 64'd89028984832, - 64'd33304588288, 64'd696442752, 64'd1099835648, - 64'd72147369984, - 64'd34130106368, - 64'd132287264, 64'd1017054656, - 64'd54991368192, - 64'd34405605376, - 64'd918431360, 64'd923245120, - 64'd37830623232, - 64'd34153697280, - 64'd1652383616, 64'd820334336, - 64'd20921751552, - 64'd33403754496, - 64'd2325779200, 64'd710291456, - 64'd4505156096, - 64'd32191121408, - 64'd2931558144, 64'd595095744, 64'd11197762560, - 64'd30556315648, - 64'd3464007424, 64'd476707168, 64'd25986973696, - 64'd28544169984, - 64'd3918779648, 64'd357038080, 64'd39685758976, - 64'd26202953728, - 64'd4292892928, 64'd237927136, 64'd52142219264, - 64'd23583496192, - 64'd4584708096, 64'd121115528, 64'd63230308352, - 64'd20738297856, - 64'd4793888256, 64'd8225954, 64'd72850481152, - 64'd17720678400, - 64'd4921340416, - 64'd99255800, 64'd80929882112, - 64'd14583931904, - 64'd4969142784, - 64'd199996272, 64'd87422132224, - 64'd11380551680, - 64'd4940455936, - 64'd292826784, 64'd92306718720, - 64'd8161475072, - 64'd4839424000, - 64'd376752768, 64'd95588089856, - 64'd4975407104, - 64'd4671066112, - 64'd450960128, 64'd97294360576, - 64'd1868203392, - 64'd4441157632, - 64'd514818656, 64'd97475715072, 64'd1117672704, - 64'd4156110592, - 64'd567882368, 64'd96202661888, 64'd3943618816, - 64'd3822844416, - 64'd609887296, 64'd93563920384, 64'd6575279616, - 64'd3448660480, - 64'd640746624, 64'd89664290816, 64'd8982853632, - 64'd3041114624, - 64'd660543296, 64'd84622270464, 64'd11141313536, - 64'd2607892992, - 64'd669520576, 64'd78567653376, 64'd13030548480, - 64'd2156690432, - 64'd668070912, 64'd71639048192, 64'd14635427840, - 64'd1695096320, - 64'd656722496, 64'd63981359104, 64'd15945781248, - 64'd1230487168, - 64'd636125120, 64'd55743389696, 64'd16956310528, - 64'd769926784, - 64'd607034560, 64'd47075373056, 64'd17666437120, - 64'd320076672, - 64'd570296128, 64'd38126714880, 64'd18080073728, 64'd112883712, - 64'd526827904, 64'd29043789824, 64'd18205360128, 64'd523325280, - 64'd477603552, 64'd19967913984, 64'd18054326272, 64'd906226560, - 64'd423635072, 64'd11033488384, 64'd17642536960, 64'd1257218688, - 64'd365956000, 64'd2366337280, 64'd16988678144, 64'd1572619008, - 64'd305604928, - 64'd5917753856, 64'd16114135040, 64'd1849452416, - 64'd243609840, - 64'd13714274304, 64'd15042542592, 64'd2085461632, - 64'd180973392, - 64'd20930994176, 64'd13799323648, 64'd2279105536, - 64'd118659216, - 64'd27488749568, 64'd12411227136, 64'd2429548288, - 64'd57579436, - 64'd33321981952, 64'd10905863168, 64'd2536636160, 64'd1416332, - 64'd38379057152, 64'd9311252480, 64'd2600868864, 64'd57550620, - 64'd42622369792, 64'd7655389184, 64'd2623358208, 64'd110126160, - 64'd46028210176, 64'd5965828096, 64'd2605783808, 64'd158532384, - 64'd48586457088, 64'd4269294080, 64'd2550340352, 64'd202250272, - 64'd50300067840, 64'd2591324928, 64'd2459678464, 64'd240855680, - 64'd51184402432, 64'd955949696, 64'd2336845568, 64'd274021024, - 64'd51266400256, - 64'd614595456, 64'd2185219584, 64'd301515488, - 64'd50583621632, - 64'd2100111616, 64'd2008443648, 64'd323203744, - 64'd49183158272, - 64'd3482639104, 64'd1810359040, 64'd339043456, - 64'd47120510976, - 64'd4746615808, 64'd1594937984, 64'd349081184, - 64'd44458311680, - 64'd5878992384, 64'd1366218752, 64'd353447680, - 64'd41265094656, - 64'd6869306880, 64'd1128242432, 64'd352351648, - 64'd37613957120, - 64'd7709711872, 64'd884992128, 64'd346072928, - 64'd33581264896, - 64'd8394967040, 64'd640337408, 64'd334954976, - 64'd29245374464, - 64'd8922391552, 64'd397981504, 64'd319396544, - 64'd24685348864, - 64'd9291779072, 64'd161414864, 64'd299843200, - 64'd19979759616, - 64'd9505280000, - 64'd66126916, 64'd276778400, - 64'd15205549056, - 64'd9567258624, - 64'd281698560, 64'd250714416, - 64'd10436952064, - 64'd9484120064, - 64'd482674976, 64'd222183376, - 64'd5744536576, - 64'd9264114688, - 64'd666774848, 64'd191728400, - 64'd1194323712, - 64'd8917130240, - 64'd832077888, 64'd159894976, 64'd3152969728, - 64'd8454461440, - 64'd977035904, 64'd127222720, 64'd7242577408, - 64'd7888576000, - 64'd1100477824, 64'd94237664, 64'd11026210816, - 64'd7232873984, - 64'd1201609088, 64'd61445076, 64'd14462461952, - 64'd6501441024, - 64'd1280004864, 64'd29322966, 64'd17517086720, - 64'd5708808704, - 64'd1335598848, - 64'd1683714, 64'd20163170304, - 64'd4869714432, - 64'd1368667008, - 64'd31168090, 64'd22381168640, - 64'd3998873344, - 64'd1379806336, - 64'd58765564, 64'd24158840832, - 64'd3110761984, - 64'd1369911040, - 64'd84157200, 64'd25491087360, - 64'd2219412736, - 64'd1340144896, - 64'd107072248, 64'd26379669504, - 64'd1338227968, - 64'd1291910528, - 64'd127289848, 64'd26832861184, - 64'd479810912, - 64'd1226817152, - 64'd144639904, 64'd26865000448, 64'd344182848, - 64'd1146647168, - 64'd159003152, 64'd26495991808, 64'd1123172992, - 64'd1053320256, - 64'd170310480, 64'd25750740992, 64'd1847759488, - 64'd948859328, - 64'd178541536, 64'd24658536448, 64'd2509805568, - 64'd835354880, - 64'd183722656, 64'd23252410368, 64'd3102496768, - 64'd714930688, - 64'd185924240, 64'd21568458752, 64'd3620379904, - 64'd589710656, - 64'd185257568, 64'd19645161472, 64'd4059376128, - 64'd461787456, - 64'd181871168, 64'd17522694144, 64'd4416777216, - 64'd333192640, - 64'd175946800, 64'd15242254336, 64'd4691217920, - 64'd205869584, - 64'd167695168, 64'd12845386752, 64'd4882632192, - 64'd81648800, - 64'd157351376, 64'd10373361664, 64'd4992191488, 64'd37773780, - 64'd145170240, 64'd7866569728, 64'd5022226432, 64'd150855536, - 64'd131421576, 64'd5363962880, 64'd4976137216, 64'd256222624, - 64'd116385472, 64'd2902548480, 64'd4858291712, 64'd352682304, - 64'd100347592, 64'd516930752, 64'd4673911808, 64'd439231904, - 64'd83594680, - 64'd1761086592, 64'd4428957184, 64'd515064448, - 64'd66410244, - 64'd3902837248, 64'd4129998080, 64'd579571264, - 64'd49070508, - 64'd5883067392, 64'd3784090880, 64'd632341440, - 64'd31840648, - 64'd7680145408, 64'd3398648064, 64'd673158400, - 64'd14971387, - 64'd9276208128, 64'd2981311488, 64'd701993600, 64'd1304030, - 64'd10657245184, 64'd2539827456, 64'd718998080, 64'd16772460, - 64'd11813120000, 64'd2081926272, 64'd724491200, 64'd31243058, - 64'd12737531904, 64'd1615208960, 64'd718948160, 64'd44549036, - 64'd13427928064, 64'd1147039616, 64'd702985152, 64'd56548972, - 64'd13885356032, 64'd684448128, 64'd677343360, 64'd67127696, - 64'd14114276352, 64'd234041408, 64'd642872064, 64'd76196728, - 64'd14122331136, - 64'd198074304, 64'd600510656, 64'd83694304, - 64'd13920076800, - 64'd606359808, 64'd551270464, 64'd89584992, - 64'd13520683008, - 64'd985897920, 64'd496216000, 64'd93858968, - 64'd12939616256, - 64'd1332436736, 64'd436446816, 64'd96530904, - 64'd12194294784, - 64'd1642420224, 64'd373079424, 64'd97638568, - 64'd11303736320, - 64'd1913007616, 64'd307229664, 64'd97241152, - 64'd10288197632, - 64'd2142081536, 64'd239996480, 64'd95417360, - 64'd9168815104, - 64'd2328243456, 64'd172446144, 64'd92263288, - 64'd7967245824, - 64'd2470800640, 64'd105598096, 64'd87890152, - 64'd6705322496, - 64'd2569741824, 64'd40412068, 64'd82421920, - 64'd5404718592, - 64'd2625704960, - 64'd22223332, 64'd75992832, - 64'd4086636288, - 64'd2639935744, - 64'd81500376, 64'd68744912, - 64'd2771511296, - 64'd2614240000, - 64'd136700320, 64'd60825504, - 64'd1478748032, - 64'd2550929664, - 64'd187199744, 64'd52384792, - 64'd226480688, - 64'd2452763904, - 64'd232475280, 64'd43573456, 64'd968635264, - 64'd2322886656, - 64'd272106496, 64'd34540396, 64'd2091598976, - 64'd2164761856, - 64'd305777152, 64'd25430600, 64'd3129207040, - 64'd1982104576, - 64'd333274944, 64'd16383198, 64'd4070163456, - 64'd1778816128, - 64'd354489568, 64'd7529658, 64'd4905154048, - 64'd1558915200, - 64'd369409440, - 64'd1007791, 64'd5626890240, - 64'd1326473344, - 64'd378117120, - 64'd9117525, 64'd6230119424, - 64'd1085551744, - 64'd380783488, - 64'd16699677, 64'd6711604224, - 64'd840141184, - 64'd377660960, - 64'd23667050, 64'd7070073344, - 64'd594106176, - 64'd369075840, - 64'd29945802, 64'd7306144768, - 64'd351133920, - 64'd355419776, - 64'd35475892, 64'd7422226432, - 64'd114687632, - 64'd337140928, - 64'd40211324, 64'd7422393344, 64'd112033768, - 64'd314734464, - 64'd44120116, 64'd7312246272, 64'd326130592, - 64'd288732960, - 64'd47184140, 64'd7098754048, 64'd525031008, - 64'd259696704, - 64'd49398688, 64'd6790086144, 64'd706513344, - 64'd228203968, - 64'd50771912, 64'd6395430400, 64'd868722176, - 64'd194841632, - 64'd51324076, 64'd5924809216, 64'd1010178368, - 64'd160195936, - 64'd51086660, 64'd5388889600, 64'd1129782656, - 64'd124843896, - 64'd50101372, 64'd4798793216, 64'd1226813696, - 64'd89345112, - 64'd48419008, 64'd4165909504, 64'd1300920576, - 64'd54234316, - 64'd46098272, 64'd3501712896, 64'd1352110080, - 64'd20014620, - 64'd43204520, 64'd2817588480, 64'd1380729216, 64'd12848429, - 64'd39808472, 64'd2124667904, 64'd1387443840, 64'd43931956, - 64'd35984880, 64'd1433674624, 64'd1373212928, 64'd72859984, - 64'd31811254, 64'd754785408, 64'd1339260800, 64'd99306744, - 64'd27366544, 64'd97505080, 64'd1287045248, 64'd122999096, - 64'd22729924, - 64'd529442272, 64'd1218225408, 64'd143718064, - 64'd17979584, - 64'd1118205056, 64'd1134626816, 64'd161299408, - 64'd13191634, - 64'd1661879040, 64'd1038206528, 64'd175633520, - 64'd8439054, - 64'd2154563328, 64'd931017408, 64'd186664304, - 64'd3790776, - 64'd2591400960, 64'd815173248, 64'd194387520, 64'd689153, - 64'd2968599296, 64'd692814272, 64'd198848272, 64'd4942285, - 64'd3283435520, 64'd566074048, 64'd200137952, 64'd8916367, - 64'd3534245632, 64'd437048064, 64'd198390720, 64'd12565821, - 64'd3720397056, 64'd307764608, 64'd193779344, 64'd15852098, - 64'd3842249728, 64'd180157664, 64'd186510832, 64'd18743908, - 64'd3901101056, 64'd56042756, 64'd176821664, 64'd21217340, - 64'd3899122432, - 64'd62904204, 64'd164972880, 64'd23255856, - 64'd3839284480, - 64'd175165168, 64'd151244992, 64'd24850182, - 64'd3725274112, - 64'd279394848, 64'd135932864, 64'd25998096, - 64'd3561405184, - 64'd374432320, 64'd119340704, 64'd26704114, - 64'd3352523520, - 64'd459309536, 64'd101776976, 64'd26979106, - 64'd3103910400, - 64'd533256096, 64'd83549712, 64'd26839824, - 64'd2821182208, - 64'd595701440, 64'd64961900, 64'd26308364, - 64'd2510190592, - 64'd646273472, 64'd46307240, 64'd25411584, - 64'd2176924160, - 64'd684794560, 64'd27866232, 64'd24180474, - 64'd1827413632, - 64'd711274816, 64'd9902631, 64'd22649494, - 64'd1467639296, - 64'd725902784, - 64'd7339646, 64'd20855898, - 64'd1103444736, - 64'd729034112, - 64'd23639200, 64'd18839040, - 64'd740456960, - 64'd721178112, - 64'd38799348, 64'd16639687, - 64'd384012864, - 64'd702982656, - 64'd52649852, 64'd14299354, - 64'd39094080, - 64'd675218176, - 64'd65048160, 64'd11859640, 64'd289729920, - 64'd638759936, - 64'd75880208, 64'd9361610, 64'd598349824, - 64'd594570112, - 64'd85060728, 64'd6845214, 64'd883155264, - 64'd543679424, - 64'd92533104, 64'd4348738, 64'd1141064448, - 64'd487168128, - 64'd98268856, 64'd1908327, 64'd1369544192, - 64'd426148000, - 64'd102266704, - 64'd442460, 64'd1566621312, - 64'd361743968, - 64'd104551240, - 64'd2673014, 64'd1730884992, - 64'd295076864, - 64'd105171344, - 64'd4755996, 64'd1861479936, - 64'd227247040, - 64'd104198272, - 64'd6667580, 64'd1958092800, - 64'd159318864, - 64'd101723504, - 64'd8387642, 64'd2020930560, - 64'd92306752, - 64'd97856440, - 64'd9899874, 64'd2050692096, - 64'd27162426, - 64'd92721856, - 64'd11191850, 64'd2048534272, 64'd35236140, - 64'd86457360, - 64'd12255013, 64'd2016032128, 64'd94094240, - 64'd79210688, - 64'd13084626, 64'd1955136000, 64'd148708208, - 64'd71137032, - 64'd13679647, 64'd1868123776, 64'd198471504, - 64'd62396380, - 64'd14042576, 64'd1757551104, 64'd242878960, - 64'd53150888, - 64'd14179239, 64'd1626200704, 64'd281529472, - 64'd43562384, - 64'd14098545, 64'd1477029504, 64'd314126912, - 64'd33789972, - 64'd13812199, 64'd1313116032, 64'd340479424, - 64'd23987790, - 64'd13334403, 64'd1137609600, 64'd360497184, - 64'd14302971, - 64'd12681513, 64'd953679040, 64'd374188960, - 64'd4873792, - 64'd11871698, 64'd764465536, 64'd381657056, 64'd4171960, - 64'd10924582, 64'd573036992, 64'd383091392, 64'd12718370, - 64'd9860880, 64'd382345600, 64'd378762368, 64'd20662552, - 64'd8702040, 64'd195190160, 64'd369012896, 64'd27915546, - 64'd7469884, 64'd14181419, 64'd354250016, 64'd34402964, - 64'd6186271, - 64'd158287360, 64'd334935488, 64'd40065392, - 64'd4872768, - 64'd320065568, 64'd311576480, 64'd44858552, - 64'd3550343, - 64'd469265472, 64'd284715680, 64'd48753232, - 64'd2239082, - 64'd604277632, 64'd254921632, 64'd51734980, - 64'd957937, - 64'd723781120, 64'd222779008, 64'd53803616, 64'd275508, - 64'd826749504, 64'd188879088, 64'd54972532, 64'd1445224, - 64'd912451840, 64'd153810704, 64'd55267860, 64'd2536908, - 64'd980448896, 64'd118151560, 64'd54727440, 64'd3538106, - 64'd1030586048, 64'd82460240, 64'd53399712, 64'd4438312, - 64'd1062981504, 64'd47268804, 64'd51342476, 64'd5229027, - 64'd1078011520, 64'd13076129, 64'd48621572, 64'd5903792, - 64'd1076292224, - 64'd19657844, 64'd45309532, 64'd6458186, - 64'd1058658880, - 64'd50517104, 64'd41484160, 64'd6889785, - 64'd1026142976, - 64'd79133616, 64'd37227136, 64'd7198112, - 64'd979947392, - 64'd105190464, 64'd32622598, 64'd7384546, - 64'd921419904, - 64'd128424112, 64'd27755788, 64'd7452206, - 64'd852026816, - 64'd148625712, 64'd22711724, 64'd7405830, - 64'd773324672, - 64'd165641600, 64'd17573944, 64'd7251620, - 64'd686933440, - 64'd179372880, 64'd12423344, 64'd6997082, - 64'd594508800, - 64'd189774240, 64'd7337101, 64'd6650849, - 64'd497716160, - 64'd196852080, 64'd2387700, 64'd6222502, - 64'd398205440, - 64'd200661888, - 64'd2357908, 64'd5722375, - 64'd297587040, - 64'd201305008, - 64'd6839042, 64'd5161374, - 64'd197410032, - 64'd198924992, - 64'd11001883, 64'd4550779, - 64'd99142048, - 64'd193703360, - 64'd14799945, 64'd3902064, - 64'd4151368, - 64'd185855120, - 64'd18194412, 64'd3226714, 64'd86308584, - 64'd175623888, - 64'd21154344, 64'd2536054, 64'd171112320, - 64'd163276960, - 64'd23656752, 64'd1841090, 64'd249272832, - 64'd149100128, - 64'd25686564, 64'd1152360, 64'd319949568, - 64'd133392576, - 64'd27236456, 64'd479799, 64'd382453888, - 64'd116461768, - 64'd28306596, - 64'd167379, 64'd436251808, - 64'd98618496, - 64'd28904270, - 64'd780780, 64'd480964704, - 64'd80172080, - 64'd29043436, - 64'd1352921, 64'd516367168, - 64'd61425856, - 64'd28744196, - 64'd1877293, 64'd542383168, - 64'd42672952, - 64'd28032188, - 64'd2348411, 64'd559079808, - 64'd24192414, - 64'd26937954, - 64'd2761848, 64'd566659456, - 64'd6245758, - 64'd25496234, - 64'd3114246, 64'd565450240, 64'd10926079, - 64'd23745258, - 64'd3403320, 64'd555894976, 64'd27105328, - 64'd21726004, - 64'd3627834, 64'd538539328, 64'd42099500, - 64'd19481452, - 64'd3787572, 64'd514018272, 64'd55743024, - 64'd17055856, - 64'd3883292, 64'd483042688, 64'd67898416, - 64'd14494022, - 64'd3916666, 64'd446385088, 64'd78456944, - 64'd11840614, - 64'd3890212, 64'd404864960, 64'd87338888, - 64'd9139497, - 64'd3807215, 64'd359334560, 64'd94493272, - 64'd6433125, - 64'd3671643, 64'd310664480, 64'd99897296, - 64'd3761978, - 64'd3488053, 64'd259729920, 64'd103555248, - 64'd1164054, - 64'd3261495, 64'd207397392, 64'd105497184, 64'd1325572, - 64'd2997414, 64'd154512336, 64'd105777200, 64'd3675132, - 64'd2701548, 64'd101887520, 64'd104471472, 64'd5856476, - 64'd2379832, 64'd50292516, 64'd101676088, 64'd7845314, - 64'd2038298, 64'd444425, 64'd97504608, 64'd9621392, - 64'd1682980, - 64'd47000308, 64'd92085560, 64'd11168599, - 64'd1319826, - 64'd91452696, 64'd85559808, 64'd12475003, - 64'd954611, - 64'd132396688, 64'd78077848, 64'd13532828, - 64'd592865, - 64'd169393344, 64'd69797112, 64'd14338368, - 64'd239796, - 64'd202083600, 64'd60879308, 64'd14891849, 64'd99768, - 64'd230189776, 64'd51487776, 64'd15197229, 64'd421433, - 64'd253515744, 64'd41785008, 64'd15261965, 64'd721283, - 64'd271945920, 64'd31930268, 64'd15096727, 64'd995915, - 64'd285443040, 64'd22077376, 64'd14715092, 64'd1242467, - 64'd294044992, 64'd12372688, 64'd14133192, 64'd1458633, - 64'd297860608, 64'd2953286, 64'd13369359, 64'd1642668, - 64'd297064512, - 64'd6054622, 64'd12443741, 64'd1793389, - 64'd291891584, - 64'd14537041, 64'd11377918, 64'd1910169, - 64'd282630240, - 64'd22393300, 64'd10194511, 64'd1992911, - 64'd269615840, - 64'd29536902, 64'd8916792, 64'd2042032, - 64'd253223232, - 64'd35896124, 64'd7568313, 64'd2058426};


endpackage
`endif

