`ifndef COEFFICIENTS_FX_SV_
`define COEFFICIENTS_FX_SV_
package Coefficients_Fx;
	localparam N = 4;
	localparam M = 4;
	localparam COEFF_BIAS = 48;
	localparam logic signed[63:0] Lfr[0:3] = {64'd260044322298584, 64'd260044322298584, 64'd250199359156856, 64'd250199359156856};
	localparam logic signed[63:0] Lfi[0:3] = {64'd63709058356239, - 64'd63709058356239, 64'd23763863612790, - 64'd23763863612790};
	localparam logic signed[63:0] Lbr[0:3] = {64'd260044322298584, 64'd260044322298584, 64'd250199359156856, 64'd250199359156856};
	localparam logic signed[63:0] Lbi[0:3] = {64'd63709058356239, - 64'd63709058356239, 64'd23763863612790, - 64'd23763863612790};
	localparam logic signed[63:0] Wfr[0:3] = {64'd2110376400288, 64'd2110376400288, - 64'd578258741790, - 64'd578258741790};
	localparam logic signed[63:0] Wfi[0:3] = {64'd408589991551, - 64'd408589991551, - 64'd1351482436250, 64'd1351482436250};
	localparam logic signed[63:0] Wbr[0:3] = {- 64'd2110376400288, - 64'd2110376400288, 64'd578258741790, 64'd578258741790};
	localparam logic signed[63:0] Wbi[0:3] = {- 64'd408589991551, 64'd408589991551, 64'd1351482436250, - 64'd1351482436250};
	localparam logic signed[63:0] Ffr[0:3][0:99] = '{
		'{64'd447026090898892, 64'd212438854663220, - 64'd118742543828233, 64'd2124069569436, 64'd533758530301235, 64'd135533022848291, - 64'd118937967428813, 64'd10703047855993, 64'd581791475334037, 64'd58223269241770, - 64'd112332143060694, 64'd17854542580099, 64'd592071790311447, - 64'd15043217072045, - 64'd99949579318250, 64'd23306691881691, 64'd567609059472628, - 64'd80473403784836, - 64'd83046631236375, 64'd26910435994395, 64'd513107491949946, - 64'd135082412638978, - 64'd63017771817475, 64'd28636321057066, 64'd434536248007739, - 64'd176786762555098, - 64'd41302914537121, 64'd28564786629008, 64'd338668554616821, - 64'd204437327937565, - 64'd19300971812962, 64'd26871111439034, 64'd232618865793307, - 64'd217795874622714, 64'd1706015050446, 64'd23806384650765, 64'd123404648130211, - 64'd217461885623591, 64'd20614854730038, 64'd19675966348113, 64'd17555435943798, - 64'd204758584317030, 64'd36547082216407, 64'd14816904712406, - 64'd79213051991507, - 64'd181588541123012, 64'd48877650159159, 64'd9575697086303, - 64'd162247347028074, - 64'd150269995034673, 64'd57246435877657, 64'd4287630382357, - 64'd228120425934556, - 64'd113365060893038, 64'd61553544592356, - 64'd741271444740, - 64'd274710326947550, - 64'd73510392031820, 64'd61940220084038, - 64'd5248911702712, - 64'd301196854566672, - 64'd33259721167799, 64'd58757822235866, - 64'd9027883505974, - 64'd307984362833831, 64'd5053872467819, 64'd52527777162492, - 64'd11932088439861, - 64'd296562061333053, 64'd39429994183574, 64'd43895643673106, - 64'd13879228597936, - 64'd269315760984741, 64'd68283322339743, 64'd33582475907727, - 64'd14849422929915, - 64'd229306420370595, 64'd90494479349139, 64'd22336513305056, - 64'd14880395954215, - 64'd180031283511389, 64'd105429486121670, 64'd10887921683993, - 64'd14059839679787, - 64'd125182888728224, 64'd112929682873037, - 64'd91124206832, - 64'd12515653555467, - 64'd68419894279291, 64'd113275504079299, - 64'd10019249073271, - 64'd10404821142049, - 64'd13161664303394, 64'd107128663692583, - 64'd18430382560606, - 64'd7901687681729, 64'd37583933958435, 64'd95458103966074, - 64'd24989355202166, - 64'd5186364118846},
		'{64'd447026090898895, 64'd212438854663220, - 64'd118742543828233, 64'd2124069569437, 64'd533758530301237, 64'd135533022848290, - 64'd118937967428813, 64'd10703047855993, 64'd581791475334039, 64'd58223269241769, - 64'd112332143060695, 64'd17854542580099, 64'd592071790311448, - 64'd15043217072045, - 64'd99949579318250, 64'd23306691881691, 64'd567609059472628, - 64'd80473403784836, - 64'd83046631236375, 64'd26910435994395, 64'd513107491949945, - 64'd135082412638978, - 64'd63017771817475, 64'd28636321057066, 64'd434536248007738, - 64'd176786762555098, - 64'd41302914537121, 64'd28564786629008, 64'd338668554616820, - 64'd204437327937565, - 64'd19300971812962, 64'd26871111439034, 64'd232618865793305, - 64'd217795874622713, 64'd1706015050446, 64'd23806384650765, 64'd123404648130209, - 64'd217461885623590, 64'd20614854730039, 64'd19675966348113, 64'd17555435943796, - 64'd204758584317030, 64'd36547082216407, 64'd14816904712405, - 64'd79213051991509, - 64'd181588541123011, 64'd48877650159160, 64'd9575697086303, - 64'd162247347028076, - 64'd150269995034672, 64'd57246435877657, 64'd4287630382357, - 64'd228120425934557, - 64'd113365060893037, 64'd61553544592356, - 64'd741271444740, - 64'd274710326947551, - 64'd73510392031820, 64'd61940220084038, - 64'd5248911702712, - 64'd301196854566673, - 64'd33259721167799, 64'd58757822235866, - 64'd9027883505974, - 64'd307984362833831, 64'd5053872467819, 64'd52527777162492, - 64'd11932088439861, - 64'd296562061333053, 64'd39429994183574, 64'd43895643673106, - 64'd13879228597936, - 64'd269315760984740, 64'd68283322339742, 64'd33582475907727, - 64'd14849422929915, - 64'd229306420370595, 64'd90494479349138, 64'd22336513305056, - 64'd14880395954215, - 64'd180031283511388, 64'd105429486121670, 64'd10887921683993, - 64'd14059839679786, - 64'd125182888728223, 64'd112929682873037, - 64'd91124206832, - 64'd12515653555467, - 64'd68419894279290, 64'd113275504079298, - 64'd10019249073271, - 64'd10404821142049, - 64'd13161664303393, 64'd107128663692583, - 64'd18430382560606, - 64'd7901687681729, 64'd37583933958436, 64'd95458103966074, - 64'd24989355202166, - 64'd5186364118846},
		'{- 64'd381499435822934, - 64'd183149749203428, 64'd86630310725113, - 64'd69190373392356, - 64'd458902695373391, - 64'd129665072389750, 64'd64049331425442, - 64'd58022328340034, - 64'd511675587650146, - 64'd84499465483901, 64'd44799412476610, - 64'd47988710248250, - 64'd543784288739743, - 64'd46845767678739, 64'd28580044483704, - 64'd39054905216160, - 64'd558793235388999, - 64'd15914185620461, 64'd15092630330722, - 64'd31171899696751, - 64'd559877165059646, 64'd9055847490855, 64'd4045912326934, - 64'd24280154551126, - 64'd549838303815003, 64'd28786786421583, - 64'd4839843942822, - 64'd18312898602776, - 64'd531127323585883, 64'd43956632171603, - 64'd11829738458406, - 64'd13198895251283, - 64'd505866896443196, 64'd55194741735207, - 64'd17172041390909, - 64'd8864735107129, - 64'd475876860632416, 64'd63079434735255, - 64'd21096770589913, - 64'd5236706101462, - 64'd442700181498718, 64'd68137079217993, - 64'd23814912933871, - 64'd2242290320462, - 64'd407629040574754, 64'd70842374507955, - 64'd25518174161999, 64'd188665902382, - 64'd371730518788098, 64'd71619582907508, - 64'd26379154908411, 64'd2123065174581, - 64'd335871455928119, 64'd70844493874180, - 64'd26551863096772, 64'd3623915347361, - 64'd300742169275819, 64'd68846933913660, - 64'd26172484519120, 64'd4749892176025, - 64'd266878800808924, 64'd65913662665606, - 64'd25360344245113, 64'd5555075015131, - 64'd234684135853854, 64'd62291520482412, - 64'd24219001447887, 64'd6088825612263, - 64'd204446797681384, 64'd58190715214252, - 64'd22837429275357, 64'd6395783347147, - 64'd176358773533097, 64'd53788155969265, - 64'd21291239547013, 64'd6515953399216, - 64'd150531269084509, 64'd49230759403064, - 64'd19643919338046, 64'd6484867285161, - 64'd127008921509744, 64'd44638669720789, - 64'd17948052959414, 64'd6333797966957, - 64'd105782427161130, 64'd40108347180554, - 64'd16246508498105, 64'd6090014277056, - 64'd86799659393969, 64'd35715491614608, - 64'd14573572996458, 64'd5777061734417, - 64'd69975366155584, 64'd31517777486311, - 64'd12956024577701, 64'd5415058931965, - 64'd55199546444852, 64'd27557385432158, - 64'd11414133423498, 64'd5021000566496},
		'{- 64'd381499435822942, - 64'd183149749203426, 64'd86630310725114, - 64'd69190373392357, - 64'd458902695373398, - 64'd129665072389749, 64'd64049331425443, - 64'd58022328340035, - 64'd511675587650152, - 64'd84499465483900, 64'd44799412476610, - 64'd47988710248250, - 64'd543784288739748, - 64'd46845767678738, 64'd28580044483704, - 64'd39054905216160, - 64'd558793235389003, - 64'd15914185620460, 64'd15092630330723, - 64'd31171899696752, - 64'd559877165059649, 64'd9055847490856, 64'd4045912326934, - 64'd24280154551126, - 64'd549838303815006, 64'd28786786421584, - 64'd4839843942821, - 64'd18312898602776, - 64'd531127323585885, 64'd43956632171603, - 64'd11829738458406, - 64'd13198895251283, - 64'd505866896443198, 64'd55194741735208, - 64'd17172041390908, - 64'd8864735107129, - 64'd475876860632417, 64'd63079434735256, - 64'd21096770589912, - 64'd5236706101462, - 64'd442700181498719, 64'd68137079217993, - 64'd23814912933871, - 64'd2242290320462, - 64'd407629040574755, 64'd70842374507956, - 64'd25518174161999, 64'd188665902382, - 64'd371730518788099, 64'd71619582907508, - 64'd26379154908411, 64'd2123065174581, - 64'd335871455928119, 64'd70844493874180, - 64'd26551863096772, 64'd3623915347361, - 64'd300742169275820, 64'd68846933913660, - 64'd26172484519120, 64'd4749892176025, - 64'd266878800808924, 64'd65913662665606, - 64'd25360344245113, 64'd5555075015131, - 64'd234684135853854, 64'd62291520482412, - 64'd24219001447887, 64'd6088825612263, - 64'd204446797681384, 64'd58190715214252, - 64'd22837429275357, 64'd6395783347147, - 64'd176358773533097, 64'd53788155969264, - 64'd21291239547013, 64'd6515953399216, - 64'd150531269084509, 64'd49230759403064, - 64'd19643919338046, 64'd6484867285161, - 64'd127008921509743, 64'd44638669720789, - 64'd17948052959414, 64'd6333797966957, - 64'd105782427161129, 64'd40108347180554, - 64'd16246508498105, 64'd6090014277056, - 64'd86799659393969, 64'd35715491614608, - 64'd14573572996458, 64'd5777061734417, - 64'd69975366155584, 64'd31517777486311, - 64'd12956024577702, 64'd5415058931965, - 64'd55199546444852, 64'd27557385432158, - 64'd11414133423498, 64'd5021000566496}};
	localparam logic signed[63:0] Ffi[0:3][0:99] = '{
		'{- 64'd533567343563437, 64'd268319199531273, 64'd40806399298483, - 64'd38617552633450, - 64'd391763233216732, 64'd295973605768580, 64'd10823330842762, - 64'd35196566838790, - 64'd241124635381047, 64'd304115619770321, - 64'd16921149543503, - 64'd30094278252985, - 64'd91083426468469, 64'd294139432460134, - 64'd41058086435045, - 64'd23761792882492, 64'd49860944995604, 64'd268339662245429, - 64'd60554639856555, - 64'd16677404110316, 64'd174537342246667, 64'd229694737316031, - 64'd74740970601041, - 64'd9316727700111, 64'd277385368107704, 64'd181631914810440, - 64'd83313864074646, - 64'd2125834056283, 64'd354619037236636, 64'd127789086059386, - 64'd86319101604800, 64'd4501375563121, 64'd404273670262553, 64'd71787257474300, - 64'd84115608763849, 64'd10240662946933, 64'd426144458395237, 64'd17025664908103, - 64'd77325160899457, 64'd14849307933993, 64'd421630520058064, - 64'd33490950346293, - 64'd66771889634250, 64'd18172185557523, 64'd393502344102755, - 64'd77286117357047, - 64'd53416011506822, 64'd20142269096978, 64'd345613178762969, - 64'd112502544078667, - 64'd38286108313483, 64'd20776061267300, 64'd282576163886429, - 64'd137949057384856, - 64'd22413958922888, 64'd20164697170800, 64'd209428881374639, - 64'd153105085656216, - 64'd6775395866267, 64'd18461638633504, 64'd131305651778233, - 64'd158086472252999, 64'd7760014389590, 64'd15867986338223, 64'd53135527076409, - 64'd153578252545104, 64'd20468438352873, 64'd12616474252706, - 64'd20619245390302, - 64'd140741374632523, 64'd30799172636449, 64'd8955184604941, - 64'd86173228075180, - 64'd121101164954702, 64'd38389558554133, 64'd5131938703205, - 64'd140569199757306, - 64'd96425637972125, 64'd43067752581663, 64'd1380189367788, - 64'd181767910603246, - 64'd68601556836605, 64'd44844351388378, - 64'd2092923542637, - 64'd208676939463808, - 64'd39515527107912, 64'd43894410608140, - 64'd5115879385566, - 64'd221122808118670, - 64'd10946424960205, 64'd40531797729240, - 64'd7559165348825, - 64'd219773347322937, 64'd15525785241805, 64'd35178071826709, - 64'd9338661000424, - 64'd206019480241986, 64'd38591205211614, 64'd28328186125272, - 64'd10416111893575},
		'{64'd533567343563435, - 64'd268319199531272, - 64'd40806399298483, 64'd38617552633450, 64'd391763233216730, - 64'd295973605768579, - 64'd10823330842762, 64'd35196566838790, 64'd241124635381044, - 64'd304115619770320, 64'd16921149543504, 64'd30094278252985, 64'd91083426468466, - 64'd294139432460134, 64'd41058086435046, 64'd23761792882492, - 64'd49860944995607, - 64'd268339662245428, 64'd60554639856555, 64'd16677404110316, - 64'd174537342246669, - 64'd229694737316030, 64'd74740970601041, 64'd9316727700110, - 64'd277385368107707, - 64'd181631914810439, 64'd83313864074646, 64'd2125834056283, - 64'd354619037236638, - 64'd127789086059385, 64'd86319101604800, - 64'd4501375563121, - 64'd404273670262554, - 64'd71787257474300, 64'd84115608763849, - 64'd10240662946933, - 64'd426144458395238, - 64'd17025664908103, 64'd77325160899457, - 64'd14849307933993, - 64'd421630520058064, 64'd33490950346293, 64'd66771889634250, - 64'd18172185557524, - 64'd393502344102754, 64'd77286117357047, 64'd53416011506822, - 64'd20142269096978, - 64'd345613178762968, 64'd112502544078667, 64'd38286108313483, - 64'd20776061267300, - 64'd282576163886428, 64'd137949057384855, 64'd22413958922888, - 64'd20164697170800, - 64'd209428881374638, 64'd153105085656216, 64'd6775395866267, - 64'd18461638633504, - 64'd131305651778232, 64'd158086472252998, - 64'd7760014389590, - 64'd15867986338223, - 64'd53135527076408, 64'd153578252545104, - 64'd20468438352873, - 64'd12616474252706, 64'd20619245390304, 64'd140741374632523, - 64'd30799172636449, - 64'd8955184604941, 64'd86173228075181, 64'd121101164954702, - 64'd38389558554133, - 64'd5131938703205, 64'd140569199757307, 64'd96425637972125, - 64'd43067752581663, - 64'd1380189367788, 64'd181767910603247, 64'd68601556836605, - 64'd44844351388378, 64'd2092923542637, 64'd208676939463809, 64'd39515527107912, - 64'd43894410608140, 64'd5115879385566, 64'd221122808118671, 64'd10946424960205, - 64'd40531797729240, 64'd7559165348825, 64'd219773347322937, - 64'd15525785241805, - 64'd35178071826709, 64'd9338661000424, 64'd206019480241986, - 64'd38591205211614, - 64'd28328186125272, 64'd10416111893575},
		'{64'd1418906945457094, - 64'd392464659842875, 64'd153449969882447, - 64'd41220299036508, 64'd1229038943134684, - 64'd364319248707501, 64'd143713503376945, - 64'd42481655525969, 64'd1053732940500831, - 64'd334785659286526, 64'd133152461584923, - 64'd42659982873121, 64'd893450353902612, - 64'd304720484157554, 64'd122139694577800, - 64'd41971395396667, 64'd748266480998832, - 64'd274816991535477, 64'd110981252952548, - 64'd40605071916859, 64'd617947321014362, - 64'd245624739051865, 64'd99923971589142, - 64'd38725032940552, 64'd502016842745322, - 64'd217568009401161, 64'd89162668944943, - 64'd36472047449026, 64'd399815327085236, - 64'd190962947708436, 64'd78846899638219, - 64'd33965605878578, 64'd310549457577359, - 64'd166033330115849, 64'd69087219393136, - 64'd31305907451388, 64'd233334856641900, - 64'd142924934035184, 64'd59960939212988, - 64'd28575820245928, 64'd167231770789332, - 64'd121718513736790, 64'd51517360285529, - 64'd25842781363707, 64'd111274598949025, - 64'd102441411360699, 64'd43782492959044, - 64'd23160612334245, 64'd64495937204794, - 64'd85077853909459, 64'd36763272498096, - 64'd20571231590821, 64'd25945783504498, - 64'd69578002120239, 64'd30451291550792, - 64'd18106251537521, - 64'd5293490319704, - 64'd55865828058739, 64'd24826074629692, - 64'd15788452505779, - 64'd30095832595756, - 64'd43845905506788, 64'd19857923697262, - 64'd13633129857659, - 64'd49283348787974, - 64'd33409201341945, 64'd15510366400756, - 64'd11649313722266, - 64'd63620803133700, - 64'd24437957679593, 64'd11742239843612, - 64'd9840863436197, - 64'd73812351748146, - 64'd16809754053264, 64'd8509443210057, - 64'd8207440779018, - 64'd80500118380676, - 64'd10400836775922, 64'd5766392253277, - 64'd6745367625675, - 64'd84264266955645, - 64'd5088799227417, 64'd3467207770480, - 64'd5448374748730, - 64'd85624266008074, - 64'd754692473764, 64'd1566668855429, - 64'd4308249257935, - 64'd85041078730737, 64'd2715359382097, 64'd20960056824, - 64'd3315388620505, - 64'd82920048313586, 64'd5428970158315, - 64'd1211760321431, - 64'd2459269414128, - 64'd79614281414177, 64'd7486665581009, - 64'd2170945581178, - 64'd1728838972406},
		'{- 64'd1418906945457094, 64'd392464659842874, - 64'd153449969882447, 64'd41220299036508, - 64'd1229038943134682, 64'd364319248707501, - 64'd143713503376945, 64'd42481655525969, - 64'd1053732940500829, 64'd334785659286525, - 64'd133152461584923, 64'd42659982873121, - 64'd893450353902610, 64'd304720484157553, - 64'd122139694577800, 64'd41971395396667, - 64'd748266480998829, 64'd274816991535476, - 64'd110981252952548, 64'd40605071916859, - 64'd617947321014359, 64'd245624739051864, - 64'd99923971589142, 64'd38725032940552, - 64'd502016842745319, 64'd217568009401160, - 64'd89162668944943, 64'd36472047449026, - 64'd399815327085234, 64'd190962947708436, - 64'd78846899638220, 64'd33965605878578, - 64'd310549457577356, 64'd166033330115849, - 64'd69087219393136, 64'd31305907451389, - 64'd233334856641898, 64'd142924934035184, - 64'd59960939212988, 64'd28575820245928, - 64'd167231770789330, 64'd121718513736789, - 64'd51517360285530, 64'd25842781363708, - 64'd111274598949023, 64'd102441411360699, - 64'd43782492959044, 64'd23160612334245, - 64'd64495937204792, 64'd85077853909459, - 64'd36763272498097, 64'd20571231590821, - 64'd25945783504497, 64'd69578002120239, - 64'd30451291550792, 64'd18106251537521, 64'd5293490319706, 64'd55865828058739, - 64'd24826074629692, 64'd15788452505779, 64'd30095832595757, 64'd43845905506787, - 64'd19857923697263, 64'd13633129857659, 64'd49283348787975, 64'd33409201341944, - 64'd15510366400756, 64'd11649313722266, 64'd63620803133701, 64'd24437957679593, - 64'd11742239843612, 64'd9840863436197, 64'd73812351748147, 64'd16809754053264, - 64'd8509443210057, 64'd8207440779018, 64'd80500118380677, 64'd10400836775922, - 64'd5766392253277, 64'd6745367625676, 64'd84264266955646, 64'd5088799227417, - 64'd3467207770480, 64'd5448374748730, 64'd85624266008075, 64'd754692473764, - 64'd1566668855429, 64'd4308249257935, 64'd85041078730737, - 64'd2715359382097, - 64'd20960056824, 64'd3315388620505, 64'd82920048313586, - 64'd5428970158315, 64'd1211760321431, 64'd2459269414128, 64'd79614281414177, - 64'd7486665581009, 64'd2170945581178, 64'd1728838972406}};
	localparam logic signed[63:0] Fbr[0:3][0:99] = '{
		'{- 64'd447026090898892, 64'd212438854663220, 64'd118742543828233, 64'd2124069569436, - 64'd533758530301235, 64'd135533022848291, 64'd118937967428813, 64'd10703047855993, - 64'd581791475334037, 64'd58223269241770, 64'd112332143060694, 64'd17854542580099, - 64'd592071790311447, - 64'd15043217072045, 64'd99949579318250, 64'd23306691881691, - 64'd567609059472628, - 64'd80473403784836, 64'd83046631236375, 64'd26910435994395, - 64'd513107491949946, - 64'd135082412638978, 64'd63017771817475, 64'd28636321057066, - 64'd434536248007739, - 64'd176786762555098, 64'd41302914537121, 64'd28564786629008, - 64'd338668554616821, - 64'd204437327937565, 64'd19300971812962, 64'd26871111439034, - 64'd232618865793307, - 64'd217795874622714, - 64'd1706015050446, 64'd23806384650765, - 64'd123404648130211, - 64'd217461885623591, - 64'd20614854730038, 64'd19675966348113, - 64'd17555435943798, - 64'd204758584317030, - 64'd36547082216407, 64'd14816904712406, 64'd79213051991507, - 64'd181588541123012, - 64'd48877650159159, 64'd9575697086303, 64'd162247347028074, - 64'd150269995034673, - 64'd57246435877657, 64'd4287630382357, 64'd228120425934556, - 64'd113365060893038, - 64'd61553544592356, - 64'd741271444740, 64'd274710326947550, - 64'd73510392031820, - 64'd61940220084038, - 64'd5248911702712, 64'd301196854566672, - 64'd33259721167799, - 64'd58757822235866, - 64'd9027883505974, 64'd307984362833831, 64'd5053872467819, - 64'd52527777162492, - 64'd11932088439861, 64'd296562061333053, 64'd39429994183574, - 64'd43895643673106, - 64'd13879228597936, 64'd269315760984741, 64'd68283322339743, - 64'd33582475907727, - 64'd14849422929915, 64'd229306420370595, 64'd90494479349139, - 64'd22336513305056, - 64'd14880395954215, 64'd180031283511389, 64'd105429486121670, - 64'd10887921683993, - 64'd14059839679787, 64'd125182888728224, 64'd112929682873037, 64'd91124206832, - 64'd12515653555467, 64'd68419894279291, 64'd113275504079299, 64'd10019249073271, - 64'd10404821142049, 64'd13161664303394, 64'd107128663692583, 64'd18430382560606, - 64'd7901687681729, - 64'd37583933958435, 64'd95458103966074, 64'd24989355202166, - 64'd5186364118846},
		'{- 64'd447026090898895, 64'd212438854663220, 64'd118742543828233, 64'd2124069569437, - 64'd533758530301237, 64'd135533022848290, 64'd118937967428813, 64'd10703047855993, - 64'd581791475334039, 64'd58223269241769, 64'd112332143060695, 64'd17854542580099, - 64'd592071790311448, - 64'd15043217072045, 64'd99949579318250, 64'd23306691881691, - 64'd567609059472628, - 64'd80473403784836, 64'd83046631236375, 64'd26910435994395, - 64'd513107491949945, - 64'd135082412638978, 64'd63017771817475, 64'd28636321057066, - 64'd434536248007738, - 64'd176786762555098, 64'd41302914537121, 64'd28564786629008, - 64'd338668554616820, - 64'd204437327937565, 64'd19300971812962, 64'd26871111439034, - 64'd232618865793305, - 64'd217795874622713, - 64'd1706015050446, 64'd23806384650765, - 64'd123404648130209, - 64'd217461885623590, - 64'd20614854730039, 64'd19675966348113, - 64'd17555435943796, - 64'd204758584317030, - 64'd36547082216407, 64'd14816904712405, 64'd79213051991509, - 64'd181588541123011, - 64'd48877650159160, 64'd9575697086303, 64'd162247347028076, - 64'd150269995034672, - 64'd57246435877657, 64'd4287630382357, 64'd228120425934557, - 64'd113365060893037, - 64'd61553544592356, - 64'd741271444740, 64'd274710326947551, - 64'd73510392031820, - 64'd61940220084038, - 64'd5248911702712, 64'd301196854566673, - 64'd33259721167799, - 64'd58757822235866, - 64'd9027883505974, 64'd307984362833831, 64'd5053872467819, - 64'd52527777162492, - 64'd11932088439861, 64'd296562061333053, 64'd39429994183574, - 64'd43895643673106, - 64'd13879228597936, 64'd269315760984740, 64'd68283322339742, - 64'd33582475907727, - 64'd14849422929915, 64'd229306420370595, 64'd90494479349138, - 64'd22336513305056, - 64'd14880395954215, 64'd180031283511388, 64'd105429486121670, - 64'd10887921683993, - 64'd14059839679786, 64'd125182888728223, 64'd112929682873037, 64'd91124206832, - 64'd12515653555467, 64'd68419894279290, 64'd113275504079298, 64'd10019249073271, - 64'd10404821142049, 64'd13161664303393, 64'd107128663692583, 64'd18430382560606, - 64'd7901687681729, - 64'd37583933958436, 64'd95458103966074, 64'd24989355202166, - 64'd5186364118846},
		'{64'd381499435822934, - 64'd183149749203428, - 64'd86630310725113, - 64'd69190373392356, 64'd458902695373391, - 64'd129665072389750, - 64'd64049331425442, - 64'd58022328340034, 64'd511675587650146, - 64'd84499465483901, - 64'd44799412476610, - 64'd47988710248250, 64'd543784288739743, - 64'd46845767678739, - 64'd28580044483704, - 64'd39054905216160, 64'd558793235388999, - 64'd15914185620461, - 64'd15092630330722, - 64'd31171899696751, 64'd559877165059646, 64'd9055847490855, - 64'd4045912326934, - 64'd24280154551126, 64'd549838303815003, 64'd28786786421583, 64'd4839843942822, - 64'd18312898602776, 64'd531127323585883, 64'd43956632171603, 64'd11829738458406, - 64'd13198895251283, 64'd505866896443196, 64'd55194741735207, 64'd17172041390909, - 64'd8864735107129, 64'd475876860632416, 64'd63079434735255, 64'd21096770589913, - 64'd5236706101462, 64'd442700181498718, 64'd68137079217993, 64'd23814912933871, - 64'd2242290320462, 64'd407629040574754, 64'd70842374507955, 64'd25518174161999, 64'd188665902382, 64'd371730518788098, 64'd71619582907508, 64'd26379154908411, 64'd2123065174581, 64'd335871455928119, 64'd70844493874180, 64'd26551863096772, 64'd3623915347361, 64'd300742169275819, 64'd68846933913660, 64'd26172484519120, 64'd4749892176025, 64'd266878800808924, 64'd65913662665606, 64'd25360344245113, 64'd5555075015131, 64'd234684135853854, 64'd62291520482412, 64'd24219001447887, 64'd6088825612263, 64'd204446797681384, 64'd58190715214252, 64'd22837429275357, 64'd6395783347147, 64'd176358773533097, 64'd53788155969265, 64'd21291239547013, 64'd6515953399216, 64'd150531269084509, 64'd49230759403064, 64'd19643919338046, 64'd6484867285161, 64'd127008921509744, 64'd44638669720789, 64'd17948052959414, 64'd6333797966957, 64'd105782427161130, 64'd40108347180554, 64'd16246508498105, 64'd6090014277056, 64'd86799659393969, 64'd35715491614608, 64'd14573572996458, 64'd5777061734417, 64'd69975366155584, 64'd31517777486311, 64'd12956024577701, 64'd5415058931965, 64'd55199546444852, 64'd27557385432158, 64'd11414133423498, 64'd5021000566496},
		'{64'd381499435822942, - 64'd183149749203426, - 64'd86630310725114, - 64'd69190373392357, 64'd458902695373398, - 64'd129665072389749, - 64'd64049331425443, - 64'd58022328340035, 64'd511675587650152, - 64'd84499465483900, - 64'd44799412476610, - 64'd47988710248250, 64'd543784288739748, - 64'd46845767678738, - 64'd28580044483704, - 64'd39054905216160, 64'd558793235389003, - 64'd15914185620460, - 64'd15092630330723, - 64'd31171899696752, 64'd559877165059649, 64'd9055847490856, - 64'd4045912326934, - 64'd24280154551126, 64'd549838303815006, 64'd28786786421584, 64'd4839843942821, - 64'd18312898602776, 64'd531127323585885, 64'd43956632171603, 64'd11829738458406, - 64'd13198895251283, 64'd505866896443198, 64'd55194741735208, 64'd17172041390908, - 64'd8864735107129, 64'd475876860632417, 64'd63079434735256, 64'd21096770589912, - 64'd5236706101462, 64'd442700181498719, 64'd68137079217993, 64'd23814912933871, - 64'd2242290320462, 64'd407629040574755, 64'd70842374507956, 64'd25518174161999, 64'd188665902382, 64'd371730518788099, 64'd71619582907508, 64'd26379154908411, 64'd2123065174581, 64'd335871455928119, 64'd70844493874180, 64'd26551863096772, 64'd3623915347361, 64'd300742169275820, 64'd68846933913660, 64'd26172484519120, 64'd4749892176025, 64'd266878800808924, 64'd65913662665606, 64'd25360344245113, 64'd5555075015131, 64'd234684135853854, 64'd62291520482412, 64'd24219001447887, 64'd6088825612263, 64'd204446797681384, 64'd58190715214252, 64'd22837429275357, 64'd6395783347147, 64'd176358773533097, 64'd53788155969264, 64'd21291239547013, 64'd6515953399216, 64'd150531269084509, 64'd49230759403064, 64'd19643919338046, 64'd6484867285161, 64'd127008921509743, 64'd44638669720789, 64'd17948052959414, 64'd6333797966957, 64'd105782427161129, 64'd40108347180554, 64'd16246508498105, 64'd6090014277056, 64'd86799659393969, 64'd35715491614608, 64'd14573572996458, 64'd5777061734417, 64'd69975366155584, 64'd31517777486311, 64'd12956024577702, 64'd5415058931965, 64'd55199546444852, 64'd27557385432158, 64'd11414133423498, 64'd5021000566496}};
	localparam logic signed[63:0] Fbi[0:3][0:99] = '{
		'{64'd533567343563437, 64'd268319199531273, - 64'd40806399298483, - 64'd38617552633450, 64'd391763233216732, 64'd295973605768580, - 64'd10823330842762, - 64'd35196566838790, 64'd241124635381047, 64'd304115619770321, 64'd16921149543503, - 64'd30094278252985, 64'd91083426468469, 64'd294139432460134, 64'd41058086435045, - 64'd23761792882492, - 64'd49860944995604, 64'd268339662245429, 64'd60554639856555, - 64'd16677404110316, - 64'd174537342246667, 64'd229694737316031, 64'd74740970601041, - 64'd9316727700111, - 64'd277385368107704, 64'd181631914810440, 64'd83313864074646, - 64'd2125834056283, - 64'd354619037236636, 64'd127789086059386, 64'd86319101604800, 64'd4501375563121, - 64'd404273670262553, 64'd71787257474300, 64'd84115608763849, 64'd10240662946933, - 64'd426144458395237, 64'd17025664908103, 64'd77325160899457, 64'd14849307933993, - 64'd421630520058064, - 64'd33490950346293, 64'd66771889634250, 64'd18172185557523, - 64'd393502344102755, - 64'd77286117357047, 64'd53416011506822, 64'd20142269096978, - 64'd345613178762969, - 64'd112502544078667, 64'd38286108313483, 64'd20776061267300, - 64'd282576163886429, - 64'd137949057384856, 64'd22413958922888, 64'd20164697170800, - 64'd209428881374639, - 64'd153105085656216, 64'd6775395866267, 64'd18461638633504, - 64'd131305651778233, - 64'd158086472252999, - 64'd7760014389590, 64'd15867986338223, - 64'd53135527076409, - 64'd153578252545104, - 64'd20468438352873, 64'd12616474252706, 64'd20619245390302, - 64'd140741374632523, - 64'd30799172636449, 64'd8955184604941, 64'd86173228075180, - 64'd121101164954702, - 64'd38389558554133, 64'd5131938703205, 64'd140569199757306, - 64'd96425637972125, - 64'd43067752581663, 64'd1380189367788, 64'd181767910603246, - 64'd68601556836605, - 64'd44844351388378, - 64'd2092923542637, 64'd208676939463808, - 64'd39515527107912, - 64'd43894410608140, - 64'd5115879385566, 64'd221122808118670, - 64'd10946424960205, - 64'd40531797729240, - 64'd7559165348825, 64'd219773347322937, 64'd15525785241805, - 64'd35178071826709, - 64'd9338661000424, 64'd206019480241986, 64'd38591205211614, - 64'd28328186125272, - 64'd10416111893575},
		'{- 64'd533567343563435, - 64'd268319199531272, 64'd40806399298483, 64'd38617552633450, - 64'd391763233216730, - 64'd295973605768579, 64'd10823330842762, 64'd35196566838790, - 64'd241124635381044, - 64'd304115619770320, - 64'd16921149543504, 64'd30094278252985, - 64'd91083426468466, - 64'd294139432460134, - 64'd41058086435046, 64'd23761792882492, 64'd49860944995607, - 64'd268339662245428, - 64'd60554639856555, 64'd16677404110316, 64'd174537342246669, - 64'd229694737316030, - 64'd74740970601041, 64'd9316727700110, 64'd277385368107707, - 64'd181631914810439, - 64'd83313864074646, 64'd2125834056283, 64'd354619037236638, - 64'd127789086059385, - 64'd86319101604800, - 64'd4501375563121, 64'd404273670262554, - 64'd71787257474300, - 64'd84115608763849, - 64'd10240662946933, 64'd426144458395238, - 64'd17025664908103, - 64'd77325160899457, - 64'd14849307933993, 64'd421630520058064, 64'd33490950346293, - 64'd66771889634250, - 64'd18172185557524, 64'd393502344102754, 64'd77286117357047, - 64'd53416011506822, - 64'd20142269096978, 64'd345613178762968, 64'd112502544078667, - 64'd38286108313483, - 64'd20776061267300, 64'd282576163886428, 64'd137949057384855, - 64'd22413958922888, - 64'd20164697170800, 64'd209428881374638, 64'd153105085656216, - 64'd6775395866267, - 64'd18461638633504, 64'd131305651778232, 64'd158086472252998, 64'd7760014389590, - 64'd15867986338223, 64'd53135527076408, 64'd153578252545104, 64'd20468438352873, - 64'd12616474252706, - 64'd20619245390304, 64'd140741374632523, 64'd30799172636449, - 64'd8955184604941, - 64'd86173228075181, 64'd121101164954702, 64'd38389558554133, - 64'd5131938703205, - 64'd140569199757307, 64'd96425637972125, 64'd43067752581663, - 64'd1380189367788, - 64'd181767910603247, 64'd68601556836605, 64'd44844351388378, 64'd2092923542637, - 64'd208676939463809, 64'd39515527107912, 64'd43894410608140, 64'd5115879385566, - 64'd221122808118671, 64'd10946424960205, 64'd40531797729240, 64'd7559165348825, - 64'd219773347322937, - 64'd15525785241805, 64'd35178071826709, 64'd9338661000424, - 64'd206019480241986, - 64'd38591205211614, 64'd28328186125272, 64'd10416111893575},
		'{- 64'd1418906945457094, - 64'd392464659842875, - 64'd153449969882447, - 64'd41220299036508, - 64'd1229038943134684, - 64'd364319248707501, - 64'd143713503376945, - 64'd42481655525969, - 64'd1053732940500831, - 64'd334785659286526, - 64'd133152461584923, - 64'd42659982873121, - 64'd893450353902612, - 64'd304720484157554, - 64'd122139694577800, - 64'd41971395396667, - 64'd748266480998832, - 64'd274816991535477, - 64'd110981252952548, - 64'd40605071916859, - 64'd617947321014362, - 64'd245624739051865, - 64'd99923971589142, - 64'd38725032940552, - 64'd502016842745322, - 64'd217568009401161, - 64'd89162668944943, - 64'd36472047449026, - 64'd399815327085236, - 64'd190962947708436, - 64'd78846899638219, - 64'd33965605878578, - 64'd310549457577359, - 64'd166033330115849, - 64'd69087219393136, - 64'd31305907451388, - 64'd233334856641900, - 64'd142924934035184, - 64'd59960939212988, - 64'd28575820245928, - 64'd167231770789332, - 64'd121718513736790, - 64'd51517360285529, - 64'd25842781363707, - 64'd111274598949025, - 64'd102441411360699, - 64'd43782492959044, - 64'd23160612334245, - 64'd64495937204794, - 64'd85077853909459, - 64'd36763272498096, - 64'd20571231590821, - 64'd25945783504498, - 64'd69578002120239, - 64'd30451291550792, - 64'd18106251537521, 64'd5293490319704, - 64'd55865828058739, - 64'd24826074629692, - 64'd15788452505779, 64'd30095832595756, - 64'd43845905506788, - 64'd19857923697262, - 64'd13633129857659, 64'd49283348787974, - 64'd33409201341945, - 64'd15510366400756, - 64'd11649313722266, 64'd63620803133700, - 64'd24437957679593, - 64'd11742239843612, - 64'd9840863436197, 64'd73812351748146, - 64'd16809754053264, - 64'd8509443210057, - 64'd8207440779018, 64'd80500118380676, - 64'd10400836775922, - 64'd5766392253277, - 64'd6745367625675, 64'd84264266955645, - 64'd5088799227417, - 64'd3467207770480, - 64'd5448374748730, 64'd85624266008074, - 64'd754692473764, - 64'd1566668855429, - 64'd4308249257935, 64'd85041078730737, 64'd2715359382097, - 64'd20960056824, - 64'd3315388620505, 64'd82920048313586, 64'd5428970158315, 64'd1211760321431, - 64'd2459269414128, 64'd79614281414177, 64'd7486665581009, 64'd2170945581178, - 64'd1728838972406},
		'{64'd1418906945457094, 64'd392464659842874, 64'd153449969882447, 64'd41220299036508, 64'd1229038943134682, 64'd364319248707501, 64'd143713503376945, 64'd42481655525969, 64'd1053732940500829, 64'd334785659286525, 64'd133152461584923, 64'd42659982873121, 64'd893450353902610, 64'd304720484157553, 64'd122139694577800, 64'd41971395396667, 64'd748266480998829, 64'd274816991535476, 64'd110981252952548, 64'd40605071916859, 64'd617947321014359, 64'd245624739051864, 64'd99923971589142, 64'd38725032940552, 64'd502016842745319, 64'd217568009401160, 64'd89162668944943, 64'd36472047449026, 64'd399815327085234, 64'd190962947708436, 64'd78846899638220, 64'd33965605878578, 64'd310549457577356, 64'd166033330115849, 64'd69087219393136, 64'd31305907451389, 64'd233334856641898, 64'd142924934035184, 64'd59960939212988, 64'd28575820245928, 64'd167231770789330, 64'd121718513736789, 64'd51517360285530, 64'd25842781363708, 64'd111274598949023, 64'd102441411360699, 64'd43782492959044, 64'd23160612334245, 64'd64495937204792, 64'd85077853909459, 64'd36763272498097, 64'd20571231590821, 64'd25945783504497, 64'd69578002120239, 64'd30451291550792, 64'd18106251537521, - 64'd5293490319706, 64'd55865828058739, 64'd24826074629692, 64'd15788452505779, - 64'd30095832595757, 64'd43845905506787, 64'd19857923697263, 64'd13633129857659, - 64'd49283348787975, 64'd33409201341944, 64'd15510366400756, 64'd11649313722266, - 64'd63620803133701, 64'd24437957679593, 64'd11742239843612, 64'd9840863436197, - 64'd73812351748147, 64'd16809754053264, 64'd8509443210057, 64'd8207440779018, - 64'd80500118380677, 64'd10400836775922, 64'd5766392253277, 64'd6745367625676, - 64'd84264266955646, 64'd5088799227417, 64'd3467207770480, 64'd5448374748730, - 64'd85624266008075, 64'd754692473764, 64'd1566668855429, 64'd4308249257935, - 64'd85041078730737, - 64'd2715359382097, 64'd20960056824, 64'd3315388620505, - 64'd82920048313586, - 64'd5428970158315, - 64'd1211760321431, 64'd2459269414128, - 64'd79614281414177, - 64'd7486665581009, - 64'd2170945581178, 64'd1728838972406}};
	localparam logic signed[63:0] hf[0:1199] = {64'd23445328887808, - 64'd609700675584, - 64'd781414694912, 64'd32420358144, 64'd22828963332096, - 64'd1792679870464, - 64'd698015809536, 64'd93131776000, 64'd21645282508800, - 64'd2877555736576, - 64'd540735307776, 64'd142618001408, 64'd19956590706688, - 64'd3813231820800, - 64'd324095016960, 64'd175894577152, 64'd17848067948544, - 64'd4559395618816, - 64'd65766854656, 64'd190096834560, 64'd15421865459712, - 64'd5088337723392, 64'd214961225728, 64'd184344248320, 64'd12790578282496, - 64'd5385808248832, 64'd498637406208, 64'd159511937024, 64'd10070498738176, - 64'd5450959945728, 64'd766943166464, 64'd117931614208, 64'd7375115780096, - 64'd5295467659264, 64'd1003777884160, 64'd63045935104, 64'd4809236152320, - 64'd4941964902400, 64'd1196091637760, - 64'd960168128, 64'd2464024363008, - 64'd4421955616768, 64'd1334444818432, - 64'd69527805952, 64'd413182361600, - 64'd3773371514880, 64'd1413289869312, - 64'd138071687168, - 64'd1289603121152, - 64'd3037959028736, 64'd1430988652544, - 64'd202289496064, - 64'd2611897434112, - 64'd2258660753408, 64'd1389590609920, - 64'd258419392512, - 64'd3542481895424, - 64'd1477150244864, 64'd1294409924608, - 64'd303436595200, - 64'd4090153402368, - 64'd731646590976, 64'd1153444872192, - 64'd335183904768, - 64'd4281524551680, - 64'd55112929280, 64'd976690872320, - 64'd352435765248, - 64'd4158039261184, 64'd526092140544, 64'd775397310464, - 64'd354898804736, - 64'd3772436185088, 64'd993073561600, 64'd561316560896, - 64'd343155539968, - 64'd3184909615104, 64'd1334763716608, 64'd345990561792, - 64'd318560075776, - 64'd2459208777728, 64'd1547815616512, 64'd140112986112, - 64'd283097006080, - 64'd1658902544384, 64'd1636073209856, - 64'd47003197440, - 64'd239215362048, - 64'd843997052928, 64'd1609688547328, - 64'd207831269376, - 64'd189649649664, - 64'd68069974016, 64'd1483967430656, - 64'd336898097152, - 64'd137240027136, 64'd623970680832, 64'd1278034313216, - 64'd430910275584, - 64'd84762025984, 64'd1197434339328, 64'd1013408006144, - 64'd488745107456, - 64'd34775007232, 64'd1628681535488, 64'd712577318912, - 64'd511319080960, 64'd10503629824, 64'd1905262460928, 64'd397657800704, - 64'd501352890368, 64'd49293500416, 64'd2025421537280, 64'd89196462080, - 64'd463056076800, 64'd80312926208, 64'd1997052444672, - 64'd194821013504, - 64'd401756422144, 64'd102806724608, 64'd1836218449920, - 64'd439723687936, - 64'd323500441600, 64'd116541661184, 64'd1565360521216, - 64'd634649903104, - 64'd234650468352, 64'd121772720128, 64'd1211326529536, - 64'd772779212800, - 64'd141501497344, 64'd119184908288, 64'd803346579456, - 64'd851313426432, - 64'd49937600512, 64'd109816037376, 64'd371078660096, - 64'd871232831488, 64'd34856198144, 64'd94966775808, - 64'd57175785472, - 64'd836861296640, 64'd108615467008, 64'd76104138752, - 64'd455999488000, - 64'd755284705280, 64'd168145059840, 64'd54764621824, - 64'd804069048320, - 64'd635668791296, 64'd211393396736, 64'd32462376960, - 64'd1085008904192, - 64'd488525201408, 64'd237455147008, 64'd10607328256, - 64'd1287876247552, - 64'd324972707840, 64'd246508945408, - 64'd9563192320, - 64'd1407283494912, - 64'd156035203072, 64'd239699853312, - 64'd27036633088, - 64'd1443189227520, 64'd7986115072, 64'd218978385920, - 64'd41059790848, - 64'd1400398807040, 64'd158038556672, 64'd186909687808, - 64'd51155476480, - 64'd1287834304512, 64'd286721146880, 64'd146466013184, - 64'd57122045952, - 64'd1117635084288, 64'd388554162176, 64'd100816445440, - 64'd59017400320, - 64'd904159952896, 64'd460112592896, 64'd53125627904, - 64'd57129889792, - 64'd662954770432, 64'd500028735488, 64'd6372370944, - 64'd51938975744, - 64'd409749815296, 64'd508876783616, - 64'd36803624960, - 64'd44068888576, - 64'd159541493760, 64'd488956690432, - 64'd74220847104, - 64'd34238554112, 64'd74198097920, 64'd443999977472, - 64'd104237334528, - 64'd23211016192, 64'd280149327872, 64'd378821279744, - 64'd125793337344, - 64'd11745245184, 64'd449591214080, 64'd298941087744, - 64'd138416570368, - 64'd552861056, 64'd576656769024, 64'd210203803648, - 64'd142193344512, 64'd9738231808, 64'd658401656832, 64'd118413475840, - 64'd137710403584, 64'd18611918848, 64'd694698967040, 64'd29006284800, - 64'd125973757952, 64'd25682835456, 64'd687983689728, - 64'd53224841216, - 64'd108311314432, 64'd30706008064, 64'd642874933248, - 64'd124342886400, - 64'd86266200064, 64'd33577543680, 64'd565709045760, - 64'd181410398208, - 64'd61488119808, 64'd34327158784, 64'd464019324928, - 64'd222562484224, - 64'd35628859392, 64'd33103777792, 64'd345996361728, - 64'd247011704832, - 64'd10247616512, 64'd30155677696, 64'd219962179584, - 64'd254991122432, 64'd13269340160, 64'd25806848000, 64'd93886406656, - 64'd247644504064, 64'd33771542528, 64'd20431253504, - 64'd25031665664, - 64'd226875015168, 64'd50387722240, 64'd14426711040, - 64'd130697568256, - 64'd195165093888, 64'd62549176320, 64'd8189863936, - 64'd218361675776, - 64'd155380285440, 64'd69993603072, 64'd2093617408, - 64'd284759916544, - 64'd110569930752, 64'd72751120384, - 64'd3531934464, - 64'd328156774400, - 64'd63776301056, 64'd71114891264, - 64'd8414319616, - 64'd348297035776, - 64'd17862291456, 64'd65599578112, - 64'd12348804096, - 64'd346278199296, 64'd24634335232, 64'd56891043840, - 64'd15203679232, - 64'd324358045696, 64'd61614284800, 64'd45791109120, - 64'd16920879104, - 64'd285714415616, 64'd91494334464, 64'd33160933376, - 64'd17512333312, - 64'd234175709184, 64'd113248165888, 64'd19866363904, - 64'd17052678144, - 64'd173940162560, 64'd126411546624, 64'd6728245248, - 64'd15669072896, - 64'd109300670464, 64'd131055050752, - 64'd5520017920, - 64'd13528996864, - 64'd44390739968, 64'd127728918528, - 64'd16265866240, - 64'd10826893312, 64'd17036284928, 64'd117385756672, - 64'd25040936960, - 64'd7770559488, 64'd71785160704, 64'd101287804928, - 64'd31533977600, - 64'd4568048640, 64'd117347885056, 64'd80905330688, - 64'd35593576448, - 64'd1415817088, 64'd151981244416, 64'd57812860928, - 64'd37221535744, 64'd1511350784, 64'd174733377536, 64'd33589395456, - 64'd36558143488, 64'd4068223488, 64'd185422594048, 64'd9727890432, - 64'd33860943872, 64'd6144569856, 64'd184574312448, - 64'd12441747456, - 64'd29478883328, 64'd7668095488, 64'd173323583488, - 64'd31812990976, - 64'd23823667200, 64'd8604938240, 64'd153292275712, - 64'd47544537088, - 64'd17340307456, 64'd8957926400, 64'd126449958912, - 64'd59083038720, - 64'd10478563328, 64'd8762915840, 64'd94968455168, - 64'd66167230464, - 64'd3666836992, 64'd8083590656, 64'd61078523904, - 64'd68815011840, 64'd2710225920, 64'd7005174272, 64'd26936915968, - 64'd67295813632, 64'd8329499136, 64'd5627514880, - 64'd5489684480, - 64'd62091300864, 64'd12941941760, 64'd4057995520, - 64'd34518839296, - 64'd53847633920, 64'd16379740160, 64'd2404689664, - 64'd58821324800, - 64'd43322970112, 64'd18558136320, 64'd770132160, - 64'd77463420928, - 64'd31333521408, 64'd19472338944, - 64'd754002112, - 64'd89922551808, - 64'd18701484032, 64'd19190188032, - 64'd2091090816, - 64'd96078036992, - 64'd6207546368, 64'd17841342464, - 64'd3182499840, - 64'd96179773440, 64'd5449682432, 64'd15604013056, - 64'd3989212416, - 64'd90798743552, 64'd15685716992, 64'd12690150400, - 64'd4492185088, - 64'd80763944960, 64'd24052670464, 64'd9330148352, - 64'd4691529216, - 64'd67090587648, 64'd30251796480, 64'd5757943296, - 64'd4604680704, - 64'd50904535040, 64'd34136342528, 64'd2197325824, - 64'd4263750144, - 64'd33367574528, 64'd35705446400, - 64'd1149855872, - 64'd3712296448, - 64'd15607789568, 64'd35090309120, - 64'd4113123328, - 64'd3001749248, 64'd1341528704, 64'd32534132736, - 64'd6560105472, - 64'd2187723776, 64'd16591755264, 64'd28367605760, - 64'd8400461824, - 64'd1326451328, 64'd29435807744, 64'd22981713920, - 64'd9587034112, - 64'd471510944, 64'd39371157504, 64'd16799712256, - 64'd10114425856, 64'd328974048, 64'd46108999680, 64'd10249914368, - 64'd10015333376, 64'd1034561984, 64'd49570344960, 64'd3740796672, - 64'd9355060224, 64'd1614068480, 64'd49870536704, - 64'd2360401920, - 64'd8224683520, 64'd2046464384, 64'd47294164992, - 64'd7744693248, - 64'd6733410304, 64'd2321107968, 64'd42262700032, - 64'd12173405184, - 64'd5000624128, 64'd2437363968, 64'd35297435648, - 64'd15485096960, - 64'd3148108288, 64'd2403686656, 64'd26980231168, - 64'd17597403136, - 64'd1292873984, 64'd2236273408, 64'd17914589184, - 64'd18504196096, 64'd459057600, 64'd1957403392, 64'd8689154048, - 64'd18268676096, 64'd2017653504, 64'd1593588736, - 64'd154424976, - 64'd17013165056, 64'd3312480000, 64'd1173659136, - 64'd8147907072, - 64'd14906490880, 64'd4294852608, 64'd726898368, - 64'd14916167680, - 64'd12149936128, 64'd4938539520, 64'd281330496, - 64'd20189716480, - 64'd8962665472, 64'd5239119360, - 64'd137757600, - 64'd23810004992, - 64'd5567526400, 64'd5212156928, - 64'd508997440, - 64'd25727895552, - 64'd2177987328, 64'd4890409984, - 64'd815784192, - 64'd25996036096, 64'd1013140992, 64'd4320324096, - 64'd1046769792, - 64'd24756170752, 64'd3842732032, 64'd3558081280, - 64'd1196009216, - 64'd22222551040, 64'd6183820288, 64'd2665468928, - 64'd1262784896, - 64'd18662825984, 64'd7949395456, 64'd1705821184, - 64'd1251149824, - 64'd14377679872, 64'd9093559296, 64'd740260416, - 64'd1169241728, - 64'd9680540672, 64'd9610226688, - 64'd175576560, - 64'd1028430144, - 64'd4878488064, 64'd9529680896, - 64'd994189760, - 64'd842360256, - 64'd255345984, 64'd8913379328, - 64'd1678149120, - 64'd625957952, 64'd3942288896, 64'd7847482880, - 64'd2201270016, - 64'd394456832, 64'd7515567104, 64'd6435587584, - 64'd2549034752, - 64'd162499888, 64'd10320179200, 64'd4791155712, - 64'd2718309376, 64'd56638868, 64'd12269389824, 64'd3030104832, - 64'd2716438784, 64'd251681216, 64'd13333505024, 64'd1263964544, - 64'd2559827968, 64'd413797600, 64'd13536129024, - 64'd406066848, - 64'd2272144640, 64'd536877568, 64'd12947745792, - 64'd1893909248, - 64'd1882277888, 64'd617618880, 64'd11677232128, - 64'd3132070144, - 64'd1422192256, 64'd655448768, 64'd9861994496, - 64'd4073722880, - 64'd924812736, 64'd652296128, 64'd7657416704, - 64'd4693409280, - 64'd422055360, 64'd612243584, 64'd5226284544, - 64'd4986456064, 64'd56896816, 64'd541089344, 64'd2728800000, - 64'd4967261696, 64'd486997696, 64'd445853024, 64'd313690464, - 64'd4666659328, 64'd848372416, 64'd334259200, - 64'd1889178880, - 64'd4128592384, 64'd1126958336, 64'd214229552, - 64'd3774414336, - 64'd3406360832, 64'd1314753152, 64'd93412432, - 64'd5264773632, - 64'd2558689792, 64'd1409694464, - 64'd21227336, - 64'd6312888320, - 64'd1645864832, 64'd1415211264, - 64'd123740512, - 64'd6901121024, - 64'd726144960, 64'd1339505536, - 64'd209436016, - 64'd7039737856, 64'd147366832, 64'd1194630016, - 64'd275028576, - 64'd6763667456, 64'd929260224, 64'd995433856, - 64'd318692288, - 64'd6128156672, 64'd1583674880, 64'd758449728, - 64'd340025568, - 64'd5203689472, 64'd2085435264, 64'd500790496, - 64'd339938592, - 64'd4070511872, 64'd2420469504, 64'd239118272, - 64'd320476352, - 64'd2813129472, 64'd2585553152, - 64'd11263037, - 64'd284593920, - 64'd1515079808, 64'd2587460864, - 64'd237151008, - 64'd235901360, - 64'd254263200, 64'd2441627136, - 64'd427997408, - 64'd178395376, 64'd900964160, 64'd2170441216, - 64'd576256960, - 64'd116194616, 64'd1894778624, 64'd1801308544, - 64'd677531584, - 64'd53293196, 64'd2685878784, 64'd1364609408, - 64'd730521408, 64'd6655250, 64'd3248457728, 64'd891683520, - 64'd736803968, 64'd60513464, 64'd3572198656, 64'd412951424, - 64'd700469952, 64'd105790296, 64'd3661387520, - 64'd43732924, - 64'd627650752, 64'd140721232, 64'd3533278720, - 64'd454425856, - 64'd525974176, 64'd164299792, 64'd3215874304, - 64'd800087168, - 64'd403987328, 64'd176262736, 64'd2745305088, - 64'd1067198784, - 64'd270581344, 64'd177034304, 64'd2162994432, - 64'd1248009600, - 64'd134451600, 64'd167636496, 64'd1512792960, - 64'd1340428288, - 64'd3620677, 64'd149573904, 64'd838246144, - 64'd1347603712, 64'd114955232, 64'd124701944, 64'd180140368, - 64'd1277245568, 64'd215681344, 64'd95087568, - 64'd425560448, - 64'd1140750976, 64'd294513728, 64'd62871340, - 64'd949306176, - 64'd952203200, 64'd349042080, 64'd30138278, - 64'd1369035008, - 64'd727312256, 64'd378471776, - 64'd1195706, - 64'd1670718080, - 64'd482364576, 64'd383515104, - 64'd29476984, - 64'd1848394624, - 64'd233239104, 64'd366207168, - 64'd53383516, - 64'd1903743232, 64'd5459444, 64'd329663904, - 64'd71968672, - 64'd1845258496, 64'd221111968, 64'd277801408, - 64'd84679440, - 64'd1687117696, 64'd403615552, 64'd215036304, - 64'd91350480, - 64'd1447830656, 64'd545719936, 64'd145986384, - 64'd92176640, - 64'd1148771840, 64'd643169216, 64'd75187936, - 64'd87667504, - 64'd812688384, 64'd694659456, 64'd6844931, - 64'd78588400, - 64'd462272224, 64'd701631680, - 64'd55379112, - 64'd65892352, - 64'd118871424, 64'd667928576, - 64'd108518560, - 64'd50647884, 64'd198599440, 64'd599346176, - 64'd150408320, - 64'd33967068, 64'd474505984, 64'd503117696, - 64'd179731040, - 64'd16937970, 64'd697073216, 64'd387363872, - 64'd196011488, - 64'd564881, 64'd858689408, 64'd260545440, - 64'd199563504, 64'd14280977, 64'd955943680, 64'd130948288, - 64'd191396832, 64'd26898452, 64'd989420288, 64'd6227536, - 64'd173093360, 64'd36780256, 64'd963284992, - 64'd106968904, - 64'd146662368, 64'd43623424, 64'd884706048, - 64'd203283504, - 64'd114385248, 64'd47327132, 64'd763159744, - 64'd278831744, - 64'd78659464, 64'd47979188, 64'd609670016, - 64'd331283296, - 64'd41850808, 64'd45833064, 64'd436032416, - 64'd359846944, - 64'd6161492, 64'd41277668, 64'd254067984, - 64'd365169088, 64'd26479866, 64'd34802248, 64'd74946664, - 64'd349159904, 64'd54502152, 64'd26958954, - 64'd91387640, - 64'd314764128, 64'd76747312, 64'd18325342, - 64'd236667376, - 64'd265694512, 64'd92497024, 64'd9469034, - 64'd354613120, - 64'd206146976, 64'd101471832, 64'd916285, - 64'd441102272, - 64'd140515312, 64'd103805208, - 64'd6874085, - 64'd494198880, - 64'd73121784, 64'd99996680, - 64'd13530434, - 64'd514055520, - 64'd7977426, 64'd90848432, - 64'd18781186, - 64'd502705856, 64'd51417016, 64'd77390752, - 64'd22460788, - 64'd463769472, 64'd102222136, 64'd60801548, - 64'd24509054, - 64'd402094368, 64'd142358800, 64'd42325120, - 64'd24964558, - 64'd323363424, 64'd170554288, 64'd23194872, - 64'd23953032, - 64'd233690992, 64'd186338080, 64'd4564007, - 64'd21671892, - 64'd139232896, 64'd189992256, - 64'd12552581, - 64'd18372148, - 64'd45831640, 64'd182463728, - 64'd27323022, - 64'd14338997, 64'd41287096, 64'd165246960, - 64'd39128472, - 64'd9872289, 64'd117753592, 64'd140246560, - 64'd47578112, - 64'd5268040, 64'd180221824, 64'd109629560, - 64'd52509720, - 64'd801917, 64'd226462704, 64'd75676936, - 64'd53977144, 64'd3284549, 64'd255384896, 64'd40642588, - 64'd52226664, 64'd6794482, 64'd266988608, 64'd6627446, - 64'd47664592, 64'd9582634, 64'd262261664, - 64'd24525796, - 64'd40818892, 64'd11558756, 64'd243029056, - 64'd51313160, - 64'd32297458, 64'd12687499, 64'd211769168, - 64'd72622888, - 64'd22745848, 64'd12985205, 64'd171410240, - 64'd87761488, - 64'd12806880, 64'd12514051, 64'd125120448, - 64'd96453440, - 64'd3084236, 64'd11374138, 64'd76104432, - 64'd98817096, 64'd5888237, 64'd9694168, 64'd27417088, - 64'd95320408, 64'd13670322, 64'd7621384, - 64'd18196422, - 64'd86720976, 64'd19931612, 64'd5311405, - 64'd58427688, - 64'd73995216, 64'd24459900, 64'd2918552, - 64'd91495096, - 64'd58261844, 64'd27162016, 64'd587176, - 64'd116195272, - 64'd40704560, 64'd28057804, - 64'd1555627, - 64'd131916592, - 64'd22498318, 64'd27268228, - 64'd3405623, - 64'd138617744, - 64'd4743168, 64'd24998842, - 64'd4885200, - 64'd136775712, 64'd11591339, 64'd21520008, - 64'd5945266, - 64'd127309288, 64'd25709012, 64'd17145312, - 64'd6565325, - 64'd111484488, 64'd37015916, 64'd12209552, - 64'd6751926, - 64'd90809376, 64'd45134976, 64'd7047641, - 64'd6535715, - 64'd66924960, 64'd49906816, 64'd1975484, - 64'd5967388, - 64'd41498968, 64'd51378136, - 64'd2726218, - 64'd5112892, - 64'd16128186, 64'd49779392, - 64'd6824629, - 64'd4048213, 64'd7745828, 64'd45494176, - 64'd10143492, - 64'd2854086, 64'd28904186, 64'd39022732, - 64'd12567793, - 64'd1610938, 64'd46398956, 64'd30942340, - 64'd14044487, - 64'd394329, 64'd59581416, 64'd21867046, - 64'd14579619, 64'd728888, 64'd68110552, 64'd12409147, - 64'd14232355, 64'd1703555, 64'd71943192, 64'd3144434, - 64'd13106544, 64'd2488240, 64'd71308104, - 64'd5417156, - 64'd11340540, 64'd3056290, 64'd66667040, - 64'd12854355, - 64'd9096031, 64'd3395945, 64'd58666224, - 64'd18850140, - 64'd6546590, 64'd3509589, 64'd48081924, - 64'd23199880, - 64'd3866646, 64'd3412269, 64'd35763800, - 64'd25812308, - 64'd1221457, 64'd3129628, 64'd22579454, - 64'd26703920, 64'd1241440, 64'd2695436, 64'd9363249, - 64'd25987774, 64'd3398958, 64'd2148887, - 64'd3128103, - 64'd23857842, 64'd5157146, 64'd1531852, - 64'd14251303, - 64'd20570246, 64'd6453776, 64'd886232, - 64'd23502344, - 64'd16422733, 64'd7258870, 64'd251566, - 64'd30531990, - 64'd11733726, 64'd7573330, - 64'd336995, - 64'd35150944, - 64'd6822198, 64'd7425958, - 64'd850280, - 64'd37325412, - 64'd1989434, 64'd6869144, - 64'd1266187, - 64'd37164228, 64'd2496474, 64'd5973642, - 64'd1570274, - 64'd34899040, 64'd6412746, 64'd4822777, - 64'd1755849, - 64'd30859434, 64'd9590306, 64'd3506502, - 64'd1823619, - 64'd25444778, 64'd11918309, 64'd2115634, - 64'd1780939, - 64'd19094822, 64'd13344914, 64'd736595, - 64'd1640764, - 64'd12260769, 64'd13874624, - 64'd553100, - 64'd1420372, - 64'd5378450, 64'd13562657, - 64'd1688413, - 64'd1139973, 64'd1155061, 64'd12506971, - 64'd2619306, - 64'd821272, 64'd7000404, 64'd10838605, - 64'd3312164, - 64'd486093, 64'd11889784, 64'd8711058, - 64'd3750148, - 64'd155118, 64'd15635430, 64'd6289390, - 64'd3932556, 64'd153179, 64'd18132676, 64'd3739718, - 64'd3873330, 64'd423375, 64'd19358022, 64'd1219631, - 64'd3598862, 64'd643693, 64'd19362732, - 64'd1129975, - 64'd3145305, 64'd806318, 64'd18262802, - 64'd3191350, - 64'd2555582, 64'd907472, 64'd16226172, - 64'd4874392, - 64'd1876292, 64'd947241, 64'd13458201, - 64'd6119158, - 64'd1154705, 64'd929205, 64'd10186395, - 64'd6896409, - 64'd435997, 64'd859896, 64'd6645324, - 64'd7206350, 64'd239119, 64'd748153, 64'd3062570, - 64'd7075816, 64'd836296, 64'd604388, - 64'd353585, - 64'd6554204, 64'd1328902, 64'd439849, - 64'd3424196, - 64'd5708510, 64'd1698806, 64'd265900, - 64'd6007069, - 64'd4617830, 64'd1936600, 64'd93355, - 64'd8001368, - 64'd3367694, 64'd2041308, - 64'd68078, - 64'd9349423, - 64'd2044582, 64'd2019633, - 64'd210254, - 64'd10035914, - 64'd730897, 64'd1884850, - 64'd326898, - 64'd10084704, 64'd499344, 64'd1655418, - 64'd413789, - 64'd9553749, 64'd1583931, 64'd1353435, - 64'd468808, - 64'd8528549, 64'd2474888, 64'd1003034, - 64'd491851, - 64'd7114641, 64'd3139850, 64'd628808, - 64'd484652, - 64'd5429680, 64'd3562420, 64'd254367, - 64'd450499, - 64'd3595570, 64'd3741589, - 64'd98915, - 64'd393910, - 64'd1731112, 64'd3690322, - 64'd412907, - 64'd320247, 64'd54482, 64'd3433492, - 64'd673446, - 64'd235337, 64'd1666896, 64'd3005323, - 64'd870764, - 64'd145095, 64'd3030674, 64'd2446552, - 64'd999632, - 64'd55173, 64'd4091727, 64'd1801485, - 64'd1059220, 64'd29330, 64'd4818380, 64'd1115126, - 64'd1052728, 64'd104112, 64'd5201045, 64'd430548, - 64'd986821, 64'd165833, 64'd5250664, - 64'd213378, - 64'd870917, 64'd212219, 64'd4996129, - 64'd783803, - 64'd716387, 64'd242085, 64'd4480926, - 64'd1255199, - 64'd535722, 64'd255301, 64'd3759262, - 64'd1610117, - 64'd341714, 64'd252699, 64'd2891956, - 64'd1839410, - 64'd146699, 64'd235934, 64'd1942340, - 64'd1941967, 64'd38108, 64'd207312, 64'd972408, - 64'd1924013, 64'd203139, 64'd169593, 64'd39406, - 64'd1798049, 64'd340867, 64'd125796, - 64'd806978, - 64'd1581546, 64'd446038, 64'd78997, - 64'd1526726, - 64'd1295473, 64'd515756, 64'd32150};
	localparam logic signed[63:0] hb[0:1199] = {64'd23445328887808, 64'd609700675584, - 64'd781414694912, - 64'd32420358144, 64'd22828963332096, 64'd1792679870464, - 64'd698015809536, - 64'd93131776000, 64'd21645282508800, 64'd2877555736576, - 64'd540735307776, - 64'd142618001408, 64'd19956590706688, 64'd3813231820800, - 64'd324095016960, - 64'd175894577152, 64'd17848067948544, 64'd4559395618816, - 64'd65766854656, - 64'd190096834560, 64'd15421865459712, 64'd5088337723392, 64'd214961225728, - 64'd184344248320, 64'd12790578282496, 64'd5385808248832, 64'd498637406208, - 64'd159511937024, 64'd10070498738176, 64'd5450959945728, 64'd766943166464, - 64'd117931614208, 64'd7375115780096, 64'd5295467659264, 64'd1003777884160, - 64'd63045935104, 64'd4809236152320, 64'd4941964902400, 64'd1196091637760, 64'd960168128, 64'd2464024363008, 64'd4421955616768, 64'd1334444818432, 64'd69527805952, 64'd413182361600, 64'd3773371514880, 64'd1413289869312, 64'd138071687168, - 64'd1289603121152, 64'd3037959028736, 64'd1430988652544, 64'd202289496064, - 64'd2611897434112, 64'd2258660753408, 64'd1389590609920, 64'd258419392512, - 64'd3542481895424, 64'd1477150244864, 64'd1294409924608, 64'd303436595200, - 64'd4090153402368, 64'd731646590976, 64'd1153444872192, 64'd335183904768, - 64'd4281524551680, 64'd55112929280, 64'd976690872320, 64'd352435765248, - 64'd4158039261184, - 64'd526092140544, 64'd775397310464, 64'd354898804736, - 64'd3772436185088, - 64'd993073561600, 64'd561316560896, 64'd343155539968, - 64'd3184909615104, - 64'd1334763716608, 64'd345990561792, 64'd318560075776, - 64'd2459208777728, - 64'd1547815616512, 64'd140112986112, 64'd283097006080, - 64'd1658902544384, - 64'd1636073209856, - 64'd47003197440, 64'd239215362048, - 64'd843997052928, - 64'd1609688547328, - 64'd207831269376, 64'd189649649664, - 64'd68069974016, - 64'd1483967430656, - 64'd336898097152, 64'd137240027136, 64'd623970680832, - 64'd1278034313216, - 64'd430910275584, 64'd84762025984, 64'd1197434339328, - 64'd1013408006144, - 64'd488745107456, 64'd34775007232, 64'd1628681535488, - 64'd712577318912, - 64'd511319080960, - 64'd10503629824, 64'd1905262460928, - 64'd397657800704, - 64'd501352890368, - 64'd49293500416, 64'd2025421537280, - 64'd89196462080, - 64'd463056076800, - 64'd80312926208, 64'd1997052444672, 64'd194821013504, - 64'd401756422144, - 64'd102806724608, 64'd1836218449920, 64'd439723687936, - 64'd323500441600, - 64'd116541661184, 64'd1565360521216, 64'd634649903104, - 64'd234650468352, - 64'd121772720128, 64'd1211326529536, 64'd772779212800, - 64'd141501497344, - 64'd119184908288, 64'd803346579456, 64'd851313426432, - 64'd49937600512, - 64'd109816037376, 64'd371078660096, 64'd871232831488, 64'd34856198144, - 64'd94966775808, - 64'd57175785472, 64'd836861296640, 64'd108615467008, - 64'd76104138752, - 64'd455999488000, 64'd755284705280, 64'd168145059840, - 64'd54764621824, - 64'd804069048320, 64'd635668791296, 64'd211393396736, - 64'd32462376960, - 64'd1085008904192, 64'd488525201408, 64'd237455147008, - 64'd10607328256, - 64'd1287876247552, 64'd324972707840, 64'd246508945408, 64'd9563192320, - 64'd1407283494912, 64'd156035203072, 64'd239699853312, 64'd27036633088, - 64'd1443189227520, - 64'd7986115072, 64'd218978385920, 64'd41059790848, - 64'd1400398807040, - 64'd158038556672, 64'd186909687808, 64'd51155476480, - 64'd1287834304512, - 64'd286721146880, 64'd146466013184, 64'd57122045952, - 64'd1117635084288, - 64'd388554162176, 64'd100816445440, 64'd59017400320, - 64'd904159952896, - 64'd460112592896, 64'd53125627904, 64'd57129889792, - 64'd662954770432, - 64'd500028735488, 64'd6372370944, 64'd51938975744, - 64'd409749815296, - 64'd508876783616, - 64'd36803624960, 64'd44068888576, - 64'd159541493760, - 64'd488956690432, - 64'd74220847104, 64'd34238554112, 64'd74198097920, - 64'd443999977472, - 64'd104237334528, 64'd23211016192, 64'd280149327872, - 64'd378821279744, - 64'd125793337344, 64'd11745245184, 64'd449591214080, - 64'd298941087744, - 64'd138416570368, 64'd552861056, 64'd576656769024, - 64'd210203803648, - 64'd142193344512, - 64'd9738231808, 64'd658401656832, - 64'd118413475840, - 64'd137710403584, - 64'd18611918848, 64'd694698967040, - 64'd29006284800, - 64'd125973757952, - 64'd25682835456, 64'd687983689728, 64'd53224841216, - 64'd108311314432, - 64'd30706008064, 64'd642874933248, 64'd124342886400, - 64'd86266200064, - 64'd33577543680, 64'd565709045760, 64'd181410398208, - 64'd61488119808, - 64'd34327158784, 64'd464019324928, 64'd222562484224, - 64'd35628859392, - 64'd33103777792, 64'd345996361728, 64'd247011704832, - 64'd10247616512, - 64'd30155677696, 64'd219962179584, 64'd254991122432, 64'd13269340160, - 64'd25806848000, 64'd93886406656, 64'd247644504064, 64'd33771542528, - 64'd20431253504, - 64'd25031665664, 64'd226875015168, 64'd50387722240, - 64'd14426711040, - 64'd130697568256, 64'd195165093888, 64'd62549176320, - 64'd8189863936, - 64'd218361675776, 64'd155380285440, 64'd69993603072, - 64'd2093617408, - 64'd284759916544, 64'd110569930752, 64'd72751120384, 64'd3531934464, - 64'd328156774400, 64'd63776301056, 64'd71114891264, 64'd8414319616, - 64'd348297035776, 64'd17862291456, 64'd65599578112, 64'd12348804096, - 64'd346278199296, - 64'd24634335232, 64'd56891043840, 64'd15203679232, - 64'd324358045696, - 64'd61614284800, 64'd45791109120, 64'd16920879104, - 64'd285714415616, - 64'd91494334464, 64'd33160933376, 64'd17512333312, - 64'd234175709184, - 64'd113248165888, 64'd19866363904, 64'd17052678144, - 64'd173940162560, - 64'd126411546624, 64'd6728245248, 64'd15669072896, - 64'd109300670464, - 64'd131055050752, - 64'd5520017920, 64'd13528996864, - 64'd44390739968, - 64'd127728918528, - 64'd16265866240, 64'd10826893312, 64'd17036284928, - 64'd117385756672, - 64'd25040936960, 64'd7770559488, 64'd71785160704, - 64'd101287804928, - 64'd31533977600, 64'd4568048640, 64'd117347885056, - 64'd80905330688, - 64'd35593576448, 64'd1415817088, 64'd151981244416, - 64'd57812860928, - 64'd37221535744, - 64'd1511350784, 64'd174733377536, - 64'd33589395456, - 64'd36558143488, - 64'd4068223488, 64'd185422594048, - 64'd9727890432, - 64'd33860943872, - 64'd6144569856, 64'd184574312448, 64'd12441747456, - 64'd29478883328, - 64'd7668095488, 64'd173323583488, 64'd31812990976, - 64'd23823667200, - 64'd8604938240, 64'd153292275712, 64'd47544537088, - 64'd17340307456, - 64'd8957926400, 64'd126449958912, 64'd59083038720, - 64'd10478563328, - 64'd8762915840, 64'd94968455168, 64'd66167230464, - 64'd3666836992, - 64'd8083590656, 64'd61078523904, 64'd68815011840, 64'd2710225920, - 64'd7005174272, 64'd26936915968, 64'd67295813632, 64'd8329499136, - 64'd5627514880, - 64'd5489684480, 64'd62091300864, 64'd12941941760, - 64'd4057995520, - 64'd34518839296, 64'd53847633920, 64'd16379740160, - 64'd2404689664, - 64'd58821324800, 64'd43322970112, 64'd18558136320, - 64'd770132160, - 64'd77463420928, 64'd31333521408, 64'd19472338944, 64'd754002112, - 64'd89922551808, 64'd18701484032, 64'd19190188032, 64'd2091090816, - 64'd96078036992, 64'd6207546368, 64'd17841342464, 64'd3182499840, - 64'd96179773440, - 64'd5449682432, 64'd15604013056, 64'd3989212416, - 64'd90798743552, - 64'd15685716992, 64'd12690150400, 64'd4492185088, - 64'd80763944960, - 64'd24052670464, 64'd9330148352, 64'd4691529216, - 64'd67090587648, - 64'd30251796480, 64'd5757943296, 64'd4604680704, - 64'd50904535040, - 64'd34136342528, 64'd2197325824, 64'd4263750144, - 64'd33367574528, - 64'd35705446400, - 64'd1149855872, 64'd3712296448, - 64'd15607789568, - 64'd35090309120, - 64'd4113123328, 64'd3001749248, 64'd1341528704, - 64'd32534132736, - 64'd6560105472, 64'd2187723776, 64'd16591755264, - 64'd28367605760, - 64'd8400461824, 64'd1326451328, 64'd29435807744, - 64'd22981713920, - 64'd9587034112, 64'd471510944, 64'd39371157504, - 64'd16799712256, - 64'd10114425856, - 64'd328974048, 64'd46108999680, - 64'd10249914368, - 64'd10015333376, - 64'd1034561984, 64'd49570344960, - 64'd3740796672, - 64'd9355060224, - 64'd1614068480, 64'd49870536704, 64'd2360401920, - 64'd8224683520, - 64'd2046464384, 64'd47294164992, 64'd7744693248, - 64'd6733410304, - 64'd2321107968, 64'd42262700032, 64'd12173405184, - 64'd5000624128, - 64'd2437363968, 64'd35297435648, 64'd15485096960, - 64'd3148108288, - 64'd2403686656, 64'd26980231168, 64'd17597403136, - 64'd1292873984, - 64'd2236273408, 64'd17914589184, 64'd18504196096, 64'd459057600, - 64'd1957403392, 64'd8689154048, 64'd18268676096, 64'd2017653504, - 64'd1593588736, - 64'd154424976, 64'd17013165056, 64'd3312480000, - 64'd1173659136, - 64'd8147907072, 64'd14906490880, 64'd4294852608, - 64'd726898368, - 64'd14916167680, 64'd12149936128, 64'd4938539520, - 64'd281330496, - 64'd20189716480, 64'd8962665472, 64'd5239119360, 64'd137757600, - 64'd23810004992, 64'd5567526400, 64'd5212156928, 64'd508997440, - 64'd25727895552, 64'd2177987328, 64'd4890409984, 64'd815784192, - 64'd25996036096, - 64'd1013140992, 64'd4320324096, 64'd1046769792, - 64'd24756170752, - 64'd3842732032, 64'd3558081280, 64'd1196009216, - 64'd22222551040, - 64'd6183820288, 64'd2665468928, 64'd1262784896, - 64'd18662825984, - 64'd7949395456, 64'd1705821184, 64'd1251149824, - 64'd14377679872, - 64'd9093559296, 64'd740260416, 64'd1169241728, - 64'd9680540672, - 64'd9610226688, - 64'd175576560, 64'd1028430144, - 64'd4878488064, - 64'd9529680896, - 64'd994189760, 64'd842360256, - 64'd255345984, - 64'd8913379328, - 64'd1678149120, 64'd625957952, 64'd3942288896, - 64'd7847482880, - 64'd2201270016, 64'd394456832, 64'd7515567104, - 64'd6435587584, - 64'd2549034752, 64'd162499888, 64'd10320179200, - 64'd4791155712, - 64'd2718309376, - 64'd56638868, 64'd12269389824, - 64'd3030104832, - 64'd2716438784, - 64'd251681216, 64'd13333505024, - 64'd1263964544, - 64'd2559827968, - 64'd413797600, 64'd13536129024, 64'd406066848, - 64'd2272144640, - 64'd536877568, 64'd12947745792, 64'd1893909248, - 64'd1882277888, - 64'd617618880, 64'd11677232128, 64'd3132070144, - 64'd1422192256, - 64'd655448768, 64'd9861994496, 64'd4073722880, - 64'd924812736, - 64'd652296128, 64'd7657416704, 64'd4693409280, - 64'd422055360, - 64'd612243584, 64'd5226284544, 64'd4986456064, 64'd56896816, - 64'd541089344, 64'd2728800000, 64'd4967261696, 64'd486997696, - 64'd445853024, 64'd313690464, 64'd4666659328, 64'd848372416, - 64'd334259200, - 64'd1889178880, 64'd4128592384, 64'd1126958336, - 64'd214229552, - 64'd3774414336, 64'd3406360832, 64'd1314753152, - 64'd93412432, - 64'd5264773632, 64'd2558689792, 64'd1409694464, 64'd21227336, - 64'd6312888320, 64'd1645864832, 64'd1415211264, 64'd123740512, - 64'd6901121024, 64'd726144960, 64'd1339505536, 64'd209436016, - 64'd7039737856, - 64'd147366832, 64'd1194630016, 64'd275028576, - 64'd6763667456, - 64'd929260224, 64'd995433856, 64'd318692288, - 64'd6128156672, - 64'd1583674880, 64'd758449728, 64'd340025568, - 64'd5203689472, - 64'd2085435264, 64'd500790496, 64'd339938592, - 64'd4070511872, - 64'd2420469504, 64'd239118272, 64'd320476352, - 64'd2813129472, - 64'd2585553152, - 64'd11263037, 64'd284593920, - 64'd1515079808, - 64'd2587460864, - 64'd237151008, 64'd235901360, - 64'd254263200, - 64'd2441627136, - 64'd427997408, 64'd178395376, 64'd900964160, - 64'd2170441216, - 64'd576256960, 64'd116194616, 64'd1894778624, - 64'd1801308544, - 64'd677531584, 64'd53293196, 64'd2685878784, - 64'd1364609408, - 64'd730521408, - 64'd6655250, 64'd3248457728, - 64'd891683520, - 64'd736803968, - 64'd60513464, 64'd3572198656, - 64'd412951424, - 64'd700469952, - 64'd105790296, 64'd3661387520, 64'd43732924, - 64'd627650752, - 64'd140721232, 64'd3533278720, 64'd454425856, - 64'd525974176, - 64'd164299792, 64'd3215874304, 64'd800087168, - 64'd403987328, - 64'd176262736, 64'd2745305088, 64'd1067198784, - 64'd270581344, - 64'd177034304, 64'd2162994432, 64'd1248009600, - 64'd134451600, - 64'd167636496, 64'd1512792960, 64'd1340428288, - 64'd3620677, - 64'd149573904, 64'd838246144, 64'd1347603712, 64'd114955232, - 64'd124701944, 64'd180140368, 64'd1277245568, 64'd215681344, - 64'd95087568, - 64'd425560448, 64'd1140750976, 64'd294513728, - 64'd62871340, - 64'd949306176, 64'd952203200, 64'd349042080, - 64'd30138278, - 64'd1369035008, 64'd727312256, 64'd378471776, 64'd1195706, - 64'd1670718080, 64'd482364576, 64'd383515104, 64'd29476984, - 64'd1848394624, 64'd233239104, 64'd366207168, 64'd53383516, - 64'd1903743232, - 64'd5459444, 64'd329663904, 64'd71968672, - 64'd1845258496, - 64'd221111968, 64'd277801408, 64'd84679440, - 64'd1687117696, - 64'd403615552, 64'd215036304, 64'd91350480, - 64'd1447830656, - 64'd545719936, 64'd145986384, 64'd92176640, - 64'd1148771840, - 64'd643169216, 64'd75187936, 64'd87667504, - 64'd812688384, - 64'd694659456, 64'd6844931, 64'd78588400, - 64'd462272224, - 64'd701631680, - 64'd55379112, 64'd65892352, - 64'd118871424, - 64'd667928576, - 64'd108518560, 64'd50647884, 64'd198599440, - 64'd599346176, - 64'd150408320, 64'd33967068, 64'd474505984, - 64'd503117696, - 64'd179731040, 64'd16937970, 64'd697073216, - 64'd387363872, - 64'd196011488, 64'd564881, 64'd858689408, - 64'd260545440, - 64'd199563504, - 64'd14280977, 64'd955943680, - 64'd130948288, - 64'd191396832, - 64'd26898452, 64'd989420288, - 64'd6227536, - 64'd173093360, - 64'd36780256, 64'd963284992, 64'd106968904, - 64'd146662368, - 64'd43623424, 64'd884706048, 64'd203283504, - 64'd114385248, - 64'd47327132, 64'd763159744, 64'd278831744, - 64'd78659464, - 64'd47979188, 64'd609670016, 64'd331283296, - 64'd41850808, - 64'd45833064, 64'd436032416, 64'd359846944, - 64'd6161492, - 64'd41277668, 64'd254067984, 64'd365169088, 64'd26479866, - 64'd34802248, 64'd74946664, 64'd349159904, 64'd54502152, - 64'd26958954, - 64'd91387640, 64'd314764128, 64'd76747312, - 64'd18325342, - 64'd236667376, 64'd265694512, 64'd92497024, - 64'd9469034, - 64'd354613120, 64'd206146976, 64'd101471832, - 64'd916285, - 64'd441102272, 64'd140515312, 64'd103805208, 64'd6874085, - 64'd494198880, 64'd73121784, 64'd99996680, 64'd13530434, - 64'd514055520, 64'd7977426, 64'd90848432, 64'd18781186, - 64'd502705856, - 64'd51417016, 64'd77390752, 64'd22460788, - 64'd463769472, - 64'd102222136, 64'd60801548, 64'd24509054, - 64'd402094368, - 64'd142358800, 64'd42325120, 64'd24964558, - 64'd323363424, - 64'd170554288, 64'd23194872, 64'd23953032, - 64'd233690992, - 64'd186338080, 64'd4564007, 64'd21671892, - 64'd139232896, - 64'd189992256, - 64'd12552581, 64'd18372148, - 64'd45831640, - 64'd182463728, - 64'd27323022, 64'd14338997, 64'd41287096, - 64'd165246960, - 64'd39128472, 64'd9872289, 64'd117753592, - 64'd140246560, - 64'd47578112, 64'd5268040, 64'd180221824, - 64'd109629560, - 64'd52509720, 64'd801917, 64'd226462704, - 64'd75676936, - 64'd53977144, - 64'd3284549, 64'd255384896, - 64'd40642588, - 64'd52226664, - 64'd6794482, 64'd266988608, - 64'd6627446, - 64'd47664592, - 64'd9582634, 64'd262261664, 64'd24525796, - 64'd40818892, - 64'd11558756, 64'd243029056, 64'd51313160, - 64'd32297458, - 64'd12687499, 64'd211769168, 64'd72622888, - 64'd22745848, - 64'd12985205, 64'd171410240, 64'd87761488, - 64'd12806880, - 64'd12514051, 64'd125120448, 64'd96453440, - 64'd3084236, - 64'd11374138, 64'd76104432, 64'd98817096, 64'd5888237, - 64'd9694168, 64'd27417088, 64'd95320408, 64'd13670322, - 64'd7621384, - 64'd18196422, 64'd86720976, 64'd19931612, - 64'd5311405, - 64'd58427688, 64'd73995216, 64'd24459900, - 64'd2918552, - 64'd91495096, 64'd58261844, 64'd27162016, - 64'd587176, - 64'd116195272, 64'd40704560, 64'd28057804, 64'd1555627, - 64'd131916592, 64'd22498318, 64'd27268228, 64'd3405623, - 64'd138617744, 64'd4743168, 64'd24998842, 64'd4885200, - 64'd136775712, - 64'd11591339, 64'd21520008, 64'd5945266, - 64'd127309288, - 64'd25709012, 64'd17145312, 64'd6565325, - 64'd111484488, - 64'd37015916, 64'd12209552, 64'd6751926, - 64'd90809376, - 64'd45134976, 64'd7047641, 64'd6535715, - 64'd66924960, - 64'd49906816, 64'd1975484, 64'd5967388, - 64'd41498968, - 64'd51378136, - 64'd2726218, 64'd5112892, - 64'd16128186, - 64'd49779392, - 64'd6824629, 64'd4048213, 64'd7745828, - 64'd45494176, - 64'd10143492, 64'd2854086, 64'd28904186, - 64'd39022732, - 64'd12567793, 64'd1610938, 64'd46398956, - 64'd30942340, - 64'd14044487, 64'd394329, 64'd59581416, - 64'd21867046, - 64'd14579619, - 64'd728888, 64'd68110552, - 64'd12409147, - 64'd14232355, - 64'd1703555, 64'd71943192, - 64'd3144434, - 64'd13106544, - 64'd2488240, 64'd71308104, 64'd5417156, - 64'd11340540, - 64'd3056290, 64'd66667040, 64'd12854355, - 64'd9096031, - 64'd3395945, 64'd58666224, 64'd18850140, - 64'd6546590, - 64'd3509589, 64'd48081924, 64'd23199880, - 64'd3866646, - 64'd3412269, 64'd35763800, 64'd25812308, - 64'd1221457, - 64'd3129628, 64'd22579454, 64'd26703920, 64'd1241440, - 64'd2695436, 64'd9363249, 64'd25987774, 64'd3398958, - 64'd2148887, - 64'd3128103, 64'd23857842, 64'd5157146, - 64'd1531852, - 64'd14251303, 64'd20570246, 64'd6453776, - 64'd886232, - 64'd23502344, 64'd16422733, 64'd7258870, - 64'd251566, - 64'd30531990, 64'd11733726, 64'd7573330, 64'd336995, - 64'd35150944, 64'd6822198, 64'd7425958, 64'd850280, - 64'd37325412, 64'd1989434, 64'd6869144, 64'd1266187, - 64'd37164228, - 64'd2496474, 64'd5973642, 64'd1570274, - 64'd34899040, - 64'd6412746, 64'd4822777, 64'd1755849, - 64'd30859434, - 64'd9590306, 64'd3506502, 64'd1823619, - 64'd25444778, - 64'd11918309, 64'd2115634, 64'd1780939, - 64'd19094822, - 64'd13344914, 64'd736595, 64'd1640764, - 64'd12260769, - 64'd13874624, - 64'd553100, 64'd1420372, - 64'd5378450, - 64'd13562657, - 64'd1688413, 64'd1139973, 64'd1155061, - 64'd12506971, - 64'd2619306, 64'd821272, 64'd7000404, - 64'd10838605, - 64'd3312164, 64'd486093, 64'd11889784, - 64'd8711058, - 64'd3750148, 64'd155118, 64'd15635430, - 64'd6289390, - 64'd3932556, - 64'd153179, 64'd18132676, - 64'd3739718, - 64'd3873330, - 64'd423375, 64'd19358022, - 64'd1219631, - 64'd3598862, - 64'd643693, 64'd19362732, 64'd1129975, - 64'd3145305, - 64'd806318, 64'd18262802, 64'd3191350, - 64'd2555582, - 64'd907472, 64'd16226172, 64'd4874392, - 64'd1876292, - 64'd947241, 64'd13458201, 64'd6119158, - 64'd1154705, - 64'd929205, 64'd10186395, 64'd6896409, - 64'd435997, - 64'd859896, 64'd6645324, 64'd7206350, 64'd239119, - 64'd748153, 64'd3062570, 64'd7075816, 64'd836296, - 64'd604388, - 64'd353585, 64'd6554204, 64'd1328902, - 64'd439849, - 64'd3424196, 64'd5708510, 64'd1698806, - 64'd265900, - 64'd6007069, 64'd4617830, 64'd1936600, - 64'd93355, - 64'd8001368, 64'd3367694, 64'd2041308, 64'd68078, - 64'd9349423, 64'd2044582, 64'd2019633, 64'd210254, - 64'd10035914, 64'd730897, 64'd1884850, 64'd326898, - 64'd10084704, - 64'd499344, 64'd1655418, 64'd413789, - 64'd9553749, - 64'd1583931, 64'd1353435, 64'd468808, - 64'd8528549, - 64'd2474888, 64'd1003034, 64'd491851, - 64'd7114641, - 64'd3139850, 64'd628808, 64'd484652, - 64'd5429680, - 64'd3562420, 64'd254367, 64'd450499, - 64'd3595570, - 64'd3741589, - 64'd98915, 64'd393910, - 64'd1731112, - 64'd3690322, - 64'd412907, 64'd320247, 64'd54482, - 64'd3433492, - 64'd673446, 64'd235337, 64'd1666896, - 64'd3005323, - 64'd870764, 64'd145095, 64'd3030674, - 64'd2446552, - 64'd999632, 64'd55173, 64'd4091727, - 64'd1801485, - 64'd1059220, - 64'd29330, 64'd4818380, - 64'd1115126, - 64'd1052728, - 64'd104112, 64'd5201045, - 64'd430548, - 64'd986821, - 64'd165833, 64'd5250664, 64'd213378, - 64'd870917, - 64'd212219, 64'd4996129, 64'd783803, - 64'd716387, - 64'd242085, 64'd4480926, 64'd1255199, - 64'd535722, - 64'd255301, 64'd3759262, 64'd1610117, - 64'd341714, - 64'd252699, 64'd2891956, 64'd1839410, - 64'd146699, - 64'd235934, 64'd1942340, 64'd1941967, 64'd38108, - 64'd207312, 64'd972408, 64'd1924013, 64'd203139, - 64'd169593, 64'd39406, 64'd1798049, 64'd340867, - 64'd125796, - 64'd806978, 64'd1581546, 64'd446038, - 64'd78997, - 64'd1526726, 64'd1295473, 64'd515756, - 64'd32150};
endpackage
`endif
