`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam N = 1;
	localparam M = 1;
	localparam COEFF_BIAS = 48;
	localparam logic signed[63:0] Lfr[0:0] = {64'd246939620925081};
	localparam logic signed[63:0] Lfi[0:0] = {64'd0};
	localparam logic signed[63:0] Lbr[0:0] = {64'd246939620925081};
	localparam logic signed[63:0] Lbi[0:0] = {64'd0};
	localparam logic signed[63:0] Wfr[0:0] = {- 64'd36844988291815};
	localparam logic signed[63:0] Wfi[0:0] = {64'd0};
	localparam logic signed[63:0] Wbr[0:0] = {64'd36844988291815};
	localparam logic signed[63:0] Wbi[0:0] = {64'd0};
	localparam logic signed[63:0] Ffr[0:0][0:19] = '{
		'{- 64'd131915342033077, - 64'd115730090598200, - 64'd101530676140075, - 64'd89073447918144, - 64'd78144649732068, - 64'd68556752034113, - 64'd60145234070172, - 64'd52765760833532, - 64'd46291706390121, - 64'd40611981077460, - 64'd35629125293769, - 64'd31257637168151, - 64'd27422505416002, - 64'd24057922204589, - 64'd21106153942605, - 64'd18516550617325, - 64'd16244676680381, - 64'd14251548568836, - 64'd12502965778025, - 64'd10968924007900}};
	localparam logic signed[63:0] Ffi[0:0][0:19] = '{
		'{64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0}};
	localparam logic signed[63:0] Fbr[0:0][0:19] = '{
		'{64'd131915342033077, 64'd115730090598200, 64'd101530676140075, 64'd89073447918144, 64'd78144649732068, 64'd68556752034113, 64'd60145234070172, 64'd52765760833532, 64'd46291706390121, 64'd40611981077460, 64'd35629125293769, 64'd31257637168151, 64'd27422505416002, 64'd24057922204589, 64'd21106153942605, 64'd18516550617325, 64'd16244676680381, 64'd14251548568836, 64'd12502965778025, 64'd10968924007900}};
	localparam logic signed[63:0] Fbi[0:0][0:19] = '{
		'{64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0}};
	localparam logic signed[63:0] hf[0:299] = {64'd17267677986816, 64'd15149033324544, 64'd13290334846976, 64'd11659686969344, 64'd10229110538240, 64'd8974057340928, 64'd7872992772096, 64'd6907022016512, 64'd6059570233344, 64'd5316095770624, 64'd4663841652736, 64'd4091615117312, 64'd3589597560832, 64'd3149174669312, 64'd2762789093376, 64'd2423810686976, 64'd2126423261184, 64'd1865523396608, 64'd1636634329088, 64'd1435828748288, 64'd1259660902400, 64'd1105107746816, 64'd969517432832, 64'd850563235840, 64'd746204037120, 64'd654649065472, 64'd574327422976, 64'd503860756480, 64'd442039959552, 64'd387804200960, 64'd340222869504, 64'd298479484928, 64'd261857771520, 64'd229729337344, 64'd201542877184, 64'd176814718976, 64'd155120582656, 64'd136088174592, 64'd119390945280, 64'd104742363136, 64'd91891081216, 64'd80616570880, 64'd70725386240, 64'd62047789056, 64'd54434881536, 64'd47756038144, 64'd41896644608, 64'd36756168704, 64'd32246398976, 64'd28289951744, 64'd24818937856, 64'd21773797376, 64'd19102277632, 64'd16758539264, 64'd14702362624, 64'd12898467840, 64'd11315900416, 64'd9927504896, 64'd8709456896, 64'd7640857088, 64'd6703367680, 64'd5880903168, 64'd5159350272, 64'd4526327808, 64'd3970973440, 64'd3483758080, 64'd3056321024, 64'd2681328128, 64'd2352344576, 64'd2063725440, 64'd1810518272, 64'd1588378112, 64'd1393493248, 64'd1222519680, 64'd1072523584, 64'd940931136, 64'd825484288, 64'd724202112, 64'd635346688, 64'd557393344, 64'd489004384, 64'd429006368, 64'd376369760, 64'd330191360, 64'd289678784, 64'd254136880, 64'd222955744, 64'd195600368, 64'd171601328, 64'd150546832, 64'd132075608, 64'd115870688, 64'd101654024, 64'd89181664, 64'd78239584, 64'd68640040, 64'd60218304, 64'd52829864, 64'd46347948, 64'd40661320, 64'd35672412, 64'd31295612, 64'd27455822, 64'd24087150, 64'd21131796, 64'd18539046, 64'd16264412, 64'd14268863, 64'd12518156, 64'd10982250, 64'd9634791, 64'd8452658, 64'd7415566, 64'd6505718, 64'd5707504, 64'd5007226, 64'd4392869, 64'd3853889, 64'd3381039, 64'd2966205, 64'd2602269, 64'd2282986, 64'd2002876, 64'd1757135, 64'd1541545, 64'd1352406, 64'd1186474, 64'd1040900, 64'd913188, 64'd801145, 64'd702849, 64'd616614, 64'd540959, 64'd474586, 64'd416357, 64'd365272, 64'd320456, 64'd281138, 64'd246644, 64'd216382, 64'd189833, 64'd166542, 64'd146108, 64'd128181, 64'd112454, 64'd98657, 64'd86552, 64'd75933, 64'd66616, 64'd58443, 64'd51272, 64'd44981, 64'd39462, 64'd34621, 64'd30373, 64'd26646, 64'd23377, 64'd20509, 64'd17992, 64'd15785, 64'd13848, 64'd12149, 64'd10658, 64'd9351, 64'd8203, 64'd7197, 64'd6314, 64'd5539, 64'd4860, 64'd4263, 64'd3740, 64'd3281, 64'd2879, 64'd2526, 64'd2216, 64'd1944, 64'd1705, 64'd1496, 64'd1313, 64'd1151, 64'd1010, 64'd886, 64'd778, 64'd682, 64'd598, 64'd525, 64'd461, 64'd404, 64'd355, 64'd311, 64'd273, 64'd239, 64'd210, 64'd184, 64'd162, 64'd142, 64'd124, 64'd109, 64'd96, 64'd84, 64'd74, 64'd65, 64'd57, 64'd50, 64'd44, 64'd38, 64'd34, 64'd29, 64'd26, 64'd23, 64'd20, 64'd17, 64'd15, 64'd13, 64'd12, 64'd10, 64'd9, 64'd8, 64'd7, 64'd6, 64'd5, 64'd5, 64'd4, 64'd4, 64'd3, 64'd3, 64'd2, 64'd2, 64'd2, 64'd2, 64'd1, 64'd1, 64'd1, 64'd1, 64'd1, 64'd1, 64'd1, 64'd1, 64'd1, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0};
	localparam logic signed[63:0] hb[0:299] = {64'd17267677986816, 64'd15149033324544, 64'd13290334846976, 64'd11659686969344, 64'd10229110538240, 64'd8974057340928, 64'd7872992772096, 64'd6907022016512, 64'd6059570233344, 64'd5316095770624, 64'd4663841652736, 64'd4091615117312, 64'd3589597560832, 64'd3149174669312, 64'd2762789093376, 64'd2423810686976, 64'd2126423261184, 64'd1865523396608, 64'd1636634329088, 64'd1435828748288, 64'd1259660902400, 64'd1105107746816, 64'd969517432832, 64'd850563235840, 64'd746204037120, 64'd654649065472, 64'd574327422976, 64'd503860756480, 64'd442039959552, 64'd387804200960, 64'd340222869504, 64'd298479484928, 64'd261857771520, 64'd229729337344, 64'd201542877184, 64'd176814718976, 64'd155120582656, 64'd136088174592, 64'd119390945280, 64'd104742363136, 64'd91891081216, 64'd80616570880, 64'd70725386240, 64'd62047789056, 64'd54434881536, 64'd47756038144, 64'd41896644608, 64'd36756168704, 64'd32246398976, 64'd28289951744, 64'd24818937856, 64'd21773797376, 64'd19102277632, 64'd16758539264, 64'd14702362624, 64'd12898467840, 64'd11315900416, 64'd9927504896, 64'd8709456896, 64'd7640857088, 64'd6703367680, 64'd5880903168, 64'd5159350272, 64'd4526327808, 64'd3970973440, 64'd3483758080, 64'd3056321024, 64'd2681328128, 64'd2352344576, 64'd2063725440, 64'd1810518272, 64'd1588378112, 64'd1393493248, 64'd1222519680, 64'd1072523584, 64'd940931136, 64'd825484288, 64'd724202112, 64'd635346688, 64'd557393344, 64'd489004384, 64'd429006368, 64'd376369760, 64'd330191360, 64'd289678784, 64'd254136880, 64'd222955744, 64'd195600368, 64'd171601328, 64'd150546832, 64'd132075608, 64'd115870688, 64'd101654024, 64'd89181664, 64'd78239584, 64'd68640040, 64'd60218304, 64'd52829864, 64'd46347948, 64'd40661320, 64'd35672412, 64'd31295612, 64'd27455822, 64'd24087150, 64'd21131796, 64'd18539046, 64'd16264412, 64'd14268863, 64'd12518156, 64'd10982250, 64'd9634791, 64'd8452658, 64'd7415566, 64'd6505718, 64'd5707504, 64'd5007226, 64'd4392869, 64'd3853889, 64'd3381039, 64'd2966205, 64'd2602269, 64'd2282986, 64'd2002876, 64'd1757135, 64'd1541545, 64'd1352406, 64'd1186474, 64'd1040900, 64'd913188, 64'd801145, 64'd702849, 64'd616614, 64'd540959, 64'd474586, 64'd416357, 64'd365272, 64'd320456, 64'd281138, 64'd246644, 64'd216382, 64'd189833, 64'd166542, 64'd146108, 64'd128181, 64'd112454, 64'd98657, 64'd86552, 64'd75933, 64'd66616, 64'd58443, 64'd51272, 64'd44981, 64'd39462, 64'd34621, 64'd30373, 64'd26646, 64'd23377, 64'd20509, 64'd17992, 64'd15785, 64'd13848, 64'd12149, 64'd10658, 64'd9351, 64'd8203, 64'd7197, 64'd6314, 64'd5539, 64'd4860, 64'd4263, 64'd3740, 64'd3281, 64'd2879, 64'd2526, 64'd2216, 64'd1944, 64'd1705, 64'd1496, 64'd1313, 64'd1151, 64'd1010, 64'd886, 64'd778, 64'd682, 64'd598, 64'd525, 64'd461, 64'd404, 64'd355, 64'd311, 64'd273, 64'd239, 64'd210, 64'd184, 64'd162, 64'd142, 64'd124, 64'd109, 64'd96, 64'd84, 64'd74, 64'd65, 64'd57, 64'd50, 64'd44, 64'd38, 64'd34, 64'd29, 64'd26, 64'd23, 64'd20, 64'd17, 64'd15, 64'd13, 64'd12, 64'd10, 64'd9, 64'd8, 64'd7, 64'd6, 64'd5, 64'd5, 64'd4, 64'd4, 64'd3, 64'd3, 64'd2, 64'd2, 64'd2, 64'd2, 64'd1, 64'd1, 64'd1, 64'd1, 64'd1, 64'd1, 64'd1, 64'd1, 64'd1, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0};
endpackage
`endif
