`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam N = 4;
	localparam real Lfr[0:3] = {0.96839535, 0.96839535, 0.94099504, 0.94099504};
	localparam real Lfi[0:3] = {0.11774739, -0.11774739, 0.0459428, -0.0459428};
	localparam real Lbr[0:3] = {0.96839535, 0.96839535, 0.94099504, 0.94099504};
	localparam real Lbi[0:3] = {0.11774739, -0.11774739, 0.0459428, -0.0459428};
	localparam real Wfr[0:3] = {-0.0005073145, -0.0005073145, 0.0001477943, 0.0001477943};
	localparam real Wfi[0:3] = {-3.5662757e-05, 3.5662757e-05, 0.00029798603, -0.00029798603};
	localparam real Wbr[0:3] = {0.0005073145, 0.0005073145, -0.0001477943, -0.0001477943};
	localparam real Wbi[0:3] = {3.5662757e-05, -3.5662757e-05, -0.00029798603, 0.00029798603};
	localparam real Ffr[0:3][0:79] = '{
		'{-12.139605, -2.8092604, 0.8107475, -0.020606074, -13.415458, -2.2923295, 0.81565076, -0.036769383, -14.43023, -1.7663188, 0.8081937, -0.051604748, -15.181462, -1.2394853, 0.78908473, -0.06495587, -15.670729, -0.7196991, 0.7591712, -0.07669605, -15.903421, -0.21434534, 0.7194201, -0.08672869, -15.888488, 0.26976246, 0.6708978, -0.09498722, -15.638121, 0.72645605, 0.6147496, -0.101434655, -15.167423, 1.1502728, 0.5521788, -0.10606273, -14.494044, 1.5365028, 0.48442578, -0.10889062, -13.637792, 1.8812228, 0.41274822, -0.10996331, -12.620233, 2.1813157, 0.33840117, -0.10934973, -11.46429, 2.4344788, 0.26261872, -0.10714051, -10.193835, 2.639218, 0.18659668, -0.10344564, -8.833287, 2.7948315, 0.11147655, -0.09839185, -7.4072256, 2.9013815, 0.03833126, -0.09211998, -5.9400115, 2.9596558, -0.031847477, -0.08478211, -4.455444, 2.9711227, -0.09815999, -0.07653885, -2.976426, 2.9378746, -0.1598076, -0.06755651, -1.524673, 2.8625672, -0.2160995, -0.05800431},
		'{-12.139605, -2.8092604, 0.8107475, -0.020606074, -13.415458, -2.2923295, 0.81565076, -0.036769383, -14.43023, -1.7663188, 0.8081937, -0.051604748, -15.181462, -1.2394853, 0.78908473, -0.06495587, -15.670729, -0.7196991, 0.7591712, -0.07669605, -15.903421, -0.21434534, 0.7194201, -0.08672869, -15.888488, 0.26976246, 0.6708978, -0.09498722, -15.638121, 0.72645605, 0.6147496, -0.101434655, -15.167423, 1.1502728, 0.5521788, -0.10606273, -14.494044, 1.5365028, 0.48442578, -0.10889062, -13.637792, 1.8812228, 0.41274822, -0.10996331, -12.620233, 2.1813157, 0.33840117, -0.10934973, -11.46429, 2.4344788, 0.26261872, -0.10714051, -10.193835, 2.639218, 0.18659668, -0.10344564, -8.833287, 2.7948315, 0.11147655, -0.09839185, -7.4072256, 2.9013815, 0.03833126, -0.09211998, -5.9400115, 2.9596558, -0.031847477, -0.08478211, -4.455444, 2.9711227, -0.09815999, -0.07653885, -2.976426, 2.9378746, -0.1598076, -0.06755651, -1.524673, 2.8625672, -0.2160995, -0.05800431},
		'{11.638412, 2.7024055, -0.71969664, 0.25664222, 12.877592, 2.2611244, -0.62268823, 0.2335727, 13.90545, 1.856806, -0.533103, 0.2117904, 14.739994, 1.4875565, -0.45060745, 0.1912724, 15.398291, 1.151498, -0.3748659, 0.1719913, 15.896471, 0.8467789, -0.30554265, 0.15391593, 16.249748, 0.5715802, -0.24230385, 0.1370118, 16.472437, 0.32412213, -0.18481918, 0.12124177, 16.577972, 0.10267011, -0.1327632, 0.10656655, 16.578936, -0.09446096, -0.08581681, 0.09294512, 16.487076, -0.26890278, -0.043668084, 0.08033521, 16.31334, -0.42223048, -0.0060134106, 0.06869361, 16.067905, -0.5559602, 0.027441842, 0.05797657, 15.760206, -0.67154723, 0.056982674, 0.048140094, 15.398962, -0.7703847, 0.08288393, 0.039140195, 14.992211, -0.853803, 0.10540992, 0.030933157, 14.547345, -0.92306876, 0.1248141, 0.023475746, 14.071136, -0.97938573, 0.14133891, 0.016725397, 13.569772, -1.0238947, 0.15521564, 0.01064037, 13.0488825, -1.057674, 0.16666435, 0.0051799035},
		'{11.638412, 2.7024055, -0.71969664, 0.25664222, 12.877592, 2.2611244, -0.62268823, 0.2335727, 13.90545, 1.856806, -0.533103, 0.2117904, 14.739994, 1.4875565, -0.45060745, 0.1912724, 15.398291, 1.151498, -0.3748659, 0.1719913, 15.896471, 0.8467789, -0.30554265, 0.15391593, 16.249748, 0.5715802, -0.24230385, 0.1370118, 16.472437, 0.32412213, -0.18481918, 0.12124177, 16.577972, 0.10267011, -0.1327632, 0.10656655, 16.578936, -0.09446096, -0.08581681, 0.09294512, 16.487076, -0.26890278, -0.043668084, 0.08033521, 16.31334, -0.42223048, -0.0060134106, 0.06869361, 16.067905, -0.5559602, 0.027441842, 0.05797657, 15.760206, -0.67154723, 0.056982674, 0.048140094, 15.398962, -0.7703847, 0.08288393, 0.039140195, 14.992211, -0.853803, 0.10540992, 0.030933157, 14.547345, -0.92306876, 0.1248141, 0.023475746, 14.071136, -0.97938573, 0.14133891, 0.016725397, 13.569772, -1.0238947, 0.15521564, 0.01064037, 13.0488825, -1.057674, 0.16666435, 0.0051799035}};
	localparam real Ffi[0:3][0:79] = '{
		'{14.093905, -3.636132, -0.25925523, 0.14280194, 12.219067, -3.8519964, -0.15559816, 0.13586244, 10.253252, -4.0001717, -0.054639798, 0.12723905, 8.23008, -4.081727, 0.04224977, 0.11714139, 6.1823936, -4.0986714, 0.13382715, 0.105790794, 4.141814, -4.0538774, 0.21898802, 0.09341655, 2.1383274, -3.9509947, 0.29677683, 0.08025208, 0.19991823, -3.794361, 0.36639377, 0.06653125, -1.647748, -3.5889034, 0.42719918, 0.052484885, -3.381596, -3.340036, 0.47871533, 0.03833751, -4.981358, -3.0535562, 0.5206256, 0.02430428, -6.4297385, -2.7355406, 0.55277145, 0.0105882585, -7.712528, -2.3922405, 0.57514715, -0.0026220253, -8.818667, -2.0299811, 0.58789253, -0.015154673, -9.740253, -1.6550634, 0.5912837, -0.02685617, -10.472513, -1.2736715, 0.58572245, -0.037592776, -11.013715, -0.8917875, 0.5717243, -0.047251556, -11.365051, -0.51511115, 0.54990524, -0.05574106, -11.53048, -0.14898933, 0.5209676, -0.062991634, -11.51653, 0.20164648, 0.48568568, -0.068955414},
		'{-14.093905, 3.636132, 0.25925523, -0.14280194, -12.219067, 3.8519964, 0.15559816, -0.13586244, -10.253252, 4.0001717, 0.054639798, -0.12723905, -8.23008, 4.081727, -0.04224977, -0.11714139, -6.1823936, 4.0986714, -0.13382715, -0.105790794, -4.141814, 4.0538774, -0.21898802, -0.09341655, -2.1383274, 3.9509947, -0.29677683, -0.08025208, -0.19991823, 3.794361, -0.36639377, -0.06653125, 1.647748, 3.5889034, -0.42719918, -0.052484885, 3.381596, 3.340036, -0.47871533, -0.03833751, 4.981358, 3.0535562, -0.5206256, -0.02430428, 6.4297385, 2.7355406, -0.55277145, -0.0105882585, 7.712528, 2.3922405, -0.57514715, 0.0026220253, 8.818667, 2.0299811, -0.58789253, 0.015154673, 9.740253, 1.6550634, -0.5912837, 0.02685617, 10.472513, 1.2736715, -0.58572245, 0.037592776, 11.013715, 0.8917875, -0.5717243, 0.047251556, 11.365051, 0.51511115, -0.54990524, 0.05574106, 11.53048, 0.14898933, -0.5209676, 0.062991634, 11.51653, -0.20164648, -0.48568568, 0.068955414},
		'{-41.919586, 6.134276, -1.1871881, 0.17252678, -38.91142, 5.896479, -1.150203, 0.17413771, -36.023823, 5.65244, -1.1109434, 0.1745937, -33.25938, 5.404225, -1.0698845, 0.17402205, -30.619717, 5.1536913, -1.0274582, 0.17254148, -28.105562, 4.902501, -0.98405546, 0.17026244, -25.716866, 4.6521325, -0.9400288, 0.16728744, -23.452885, 4.403894, -0.89569455, 0.16371135, -21.31226, 4.158933, -0.8513352, 0.15962176, -19.29309, 3.9182527, -0.80720174, 0.15509926, -17.39302, 3.6827166, -0.76351553, 0.15021779, -15.609284, 3.453064, -0.72047055, 0.14504503, -13.938779, 3.2299175, -0.67823553, 0.13964263, -12.378118, 3.0137942, -0.6369555, 0.13406663, -10.923679, 2.8051126, -0.596754, 0.12836772, -9.571656, 2.6042035, -0.55773467, 0.1225916, -8.318097, 2.4113164, -0.51998276, 0.11677924, -7.1589427, 2.2266283, -0.48356685, 0.11096723, -6.090062, 2.0502505, -0.4485405, 0.10518803, -5.107285, 1.882235, -0.41494337, 0.09947026},
		'{41.919586, -6.134276, 1.1871881, -0.17252678, 38.91142, -5.896479, 1.150203, -0.17413771, 36.023823, -5.65244, 1.1109434, -0.1745937, 33.25938, -5.404225, 1.0698845, -0.17402205, 30.619717, -5.1536913, 1.0274582, -0.17254148, 28.105562, -4.902501, 0.98405546, -0.17026244, 25.716866, -4.6521325, 0.9400288, -0.16728744, 23.452885, -4.403894, 0.89569455, -0.16371135, 21.31226, -4.158933, 0.8513352, -0.15962176, 19.29309, -3.9182527, 0.80720174, -0.15509926, 17.39302, -3.6827166, 0.76351553, -0.15021779, 15.609284, -3.453064, 0.72047055, -0.14504503, 13.938779, -3.2299175, 0.67823553, -0.13964263, 12.378118, -3.0137942, 0.6369555, -0.13406663, 10.923679, -2.8051126, 0.596754, -0.12836772, 9.571656, -2.6042035, 0.55773467, -0.1225916, 8.318097, -2.4113164, 0.51998276, -0.11677924, 7.1589427, -2.2266283, 0.48356685, -0.11096723, 6.090062, -2.0502505, 0.4485405, -0.10518803, 5.107285, -1.882235, 0.41494337, -0.09947026}};
	localparam real Fbr[0:3][0:79] = '{
		'{12.139605, -2.8092604, -0.8107475, -0.020606074, 13.415458, -2.2923295, -0.81565076, -0.036769383, 14.43023, -1.7663188, -0.8081937, -0.051604748, 15.181462, -1.2394853, -0.78908473, -0.06495587, 15.670729, -0.7196991, -0.7591712, -0.07669605, 15.903421, -0.21434534, -0.7194201, -0.08672869, 15.888488, 0.26976246, -0.6708978, -0.09498722, 15.638121, 0.72645605, -0.6147496, -0.101434655, 15.167423, 1.1502728, -0.5521788, -0.10606273, 14.494044, 1.5365028, -0.48442578, -0.10889062, 13.637792, 1.8812228, -0.41274822, -0.10996331, 12.620233, 2.1813157, -0.33840117, -0.10934973, 11.46429, 2.4344788, -0.26261872, -0.10714051, 10.193835, 2.639218, -0.18659668, -0.10344564, 8.833287, 2.7948315, -0.11147655, -0.09839185, 7.4072256, 2.9013815, -0.03833126, -0.09211998, 5.9400115, 2.9596558, 0.031847477, -0.08478211, 4.455444, 2.9711227, 0.09815999, -0.07653885, 2.976426, 2.9378746, 0.1598076, -0.06755651, 1.524673, 2.8625672, 0.2160995, -0.05800431},
		'{12.139605, -2.8092604, -0.8107475, -0.020606074, 13.415458, -2.2923295, -0.81565076, -0.036769383, 14.43023, -1.7663188, -0.8081937, -0.051604748, 15.181462, -1.2394853, -0.78908473, -0.06495587, 15.670729, -0.7196991, -0.7591712, -0.07669605, 15.903421, -0.21434534, -0.7194201, -0.08672869, 15.888488, 0.26976246, -0.6708978, -0.09498722, 15.638121, 0.72645605, -0.6147496, -0.101434655, 15.167423, 1.1502728, -0.5521788, -0.10606273, 14.494044, 1.5365028, -0.48442578, -0.10889062, 13.637792, 1.8812228, -0.41274822, -0.10996331, 12.620233, 2.1813157, -0.33840117, -0.10934973, 11.46429, 2.4344788, -0.26261872, -0.10714051, 10.193835, 2.639218, -0.18659668, -0.10344564, 8.833287, 2.7948315, -0.11147655, -0.09839185, 7.4072256, 2.9013815, -0.03833126, -0.09211998, 5.9400115, 2.9596558, 0.031847477, -0.08478211, 4.455444, 2.9711227, 0.09815999, -0.07653885, 2.976426, 2.9378746, 0.1598076, -0.06755651, 1.524673, 2.8625672, 0.2160995, -0.05800431},
		'{-11.638412, 2.7024055, 0.71969664, 0.25664222, -12.877592, 2.2611244, 0.62268823, 0.2335727, -13.90545, 1.856806, 0.533103, 0.2117904, -14.739994, 1.4875565, 0.45060745, 0.1912724, -15.398291, 1.151498, 0.3748659, 0.1719913, -15.896471, 0.8467789, 0.30554265, 0.15391593, -16.249748, 0.5715802, 0.24230385, 0.1370118, -16.472437, 0.32412213, 0.18481918, 0.12124177, -16.577972, 0.10267011, 0.1327632, 0.10656655, -16.578936, -0.09446096, 0.08581681, 0.09294512, -16.487076, -0.26890278, 0.043668084, 0.08033521, -16.31334, -0.42223048, 0.0060134106, 0.06869361, -16.067905, -0.5559602, -0.027441842, 0.05797657, -15.760206, -0.67154723, -0.056982674, 0.048140094, -15.398962, -0.7703847, -0.08288393, 0.039140195, -14.992211, -0.853803, -0.10540992, 0.030933157, -14.547345, -0.92306876, -0.1248141, 0.023475746, -14.071136, -0.97938573, -0.14133891, 0.016725397, -13.569772, -1.0238947, -0.15521564, 0.01064037, -13.0488825, -1.057674, -0.16666435, 0.0051799035},
		'{-11.638412, 2.7024055, 0.71969664, 0.25664222, -12.877592, 2.2611244, 0.62268823, 0.2335727, -13.90545, 1.856806, 0.533103, 0.2117904, -14.739994, 1.4875565, 0.45060745, 0.1912724, -15.398291, 1.151498, 0.3748659, 0.1719913, -15.896471, 0.8467789, 0.30554265, 0.15391593, -16.249748, 0.5715802, 0.24230385, 0.1370118, -16.472437, 0.32412213, 0.18481918, 0.12124177, -16.577972, 0.10267011, 0.1327632, 0.10656655, -16.578936, -0.09446096, 0.08581681, 0.09294512, -16.487076, -0.26890278, 0.043668084, 0.08033521, -16.31334, -0.42223048, 0.0060134106, 0.06869361, -16.067905, -0.5559602, -0.027441842, 0.05797657, -15.760206, -0.67154723, -0.056982674, 0.048140094, -15.398962, -0.7703847, -0.08288393, 0.039140195, -14.992211, -0.853803, -0.10540992, 0.030933157, -14.547345, -0.92306876, -0.1248141, 0.023475746, -14.071136, -0.97938573, -0.14133891, 0.016725397, -13.569772, -1.0238947, -0.15521564, 0.01064037, -13.0488825, -1.057674, -0.16666435, 0.0051799035}};
	localparam real Fbi[0:3][0:79] = '{
		'{-14.093905, -3.636132, 0.25925523, 0.14280194, -12.219067, -3.8519964, 0.15559816, 0.13586244, -10.253252, -4.0001717, 0.054639798, 0.12723905, -8.23008, -4.081727, -0.04224977, 0.11714139, -6.1823936, -4.0986714, -0.13382715, 0.105790794, -4.141814, -4.0538774, -0.21898802, 0.09341655, -2.1383274, -3.9509947, -0.29677683, 0.08025208, -0.19991823, -3.794361, -0.36639377, 0.06653125, 1.647748, -3.5889034, -0.42719918, 0.052484885, 3.381596, -3.340036, -0.47871533, 0.03833751, 4.981358, -3.0535562, -0.5206256, 0.02430428, 6.4297385, -2.7355406, -0.55277145, 0.0105882585, 7.712528, -2.3922405, -0.57514715, -0.0026220253, 8.818667, -2.0299811, -0.58789253, -0.015154673, 9.740253, -1.6550634, -0.5912837, -0.02685617, 10.472513, -1.2736715, -0.58572245, -0.037592776, 11.013715, -0.8917875, -0.5717243, -0.047251556, 11.365051, -0.51511115, -0.54990524, -0.05574106, 11.53048, -0.14898933, -0.5209676, -0.062991634, 11.51653, 0.20164648, -0.48568568, -0.068955414},
		'{14.093905, 3.636132, -0.25925523, -0.14280194, 12.219067, 3.8519964, -0.15559816, -0.13586244, 10.253252, 4.0001717, -0.054639798, -0.12723905, 8.23008, 4.081727, 0.04224977, -0.11714139, 6.1823936, 4.0986714, 0.13382715, -0.105790794, 4.141814, 4.0538774, 0.21898802, -0.09341655, 2.1383274, 3.9509947, 0.29677683, -0.08025208, 0.19991823, 3.794361, 0.36639377, -0.06653125, -1.647748, 3.5889034, 0.42719918, -0.052484885, -3.381596, 3.340036, 0.47871533, -0.03833751, -4.981358, 3.0535562, 0.5206256, -0.02430428, -6.4297385, 2.7355406, 0.55277145, -0.0105882585, -7.712528, 2.3922405, 0.57514715, 0.0026220253, -8.818667, 2.0299811, 0.58789253, 0.015154673, -9.740253, 1.6550634, 0.5912837, 0.02685617, -10.472513, 1.2736715, 0.58572245, 0.037592776, -11.013715, 0.8917875, 0.5717243, 0.047251556, -11.365051, 0.51511115, 0.54990524, 0.05574106, -11.53048, 0.14898933, 0.5209676, 0.062991634, -11.51653, -0.20164648, 0.48568568, 0.068955414},
		'{41.919586, 6.134276, 1.1871881, 0.17252678, 38.91142, 5.896479, 1.150203, 0.17413771, 36.023823, 5.65244, 1.1109434, 0.1745937, 33.25938, 5.404225, 1.0698845, 0.17402205, 30.619717, 5.1536913, 1.0274582, 0.17254148, 28.105562, 4.902501, 0.98405546, 0.17026244, 25.716866, 4.6521325, 0.9400288, 0.16728744, 23.452885, 4.403894, 0.89569455, 0.16371135, 21.31226, 4.158933, 0.8513352, 0.15962176, 19.29309, 3.9182527, 0.80720174, 0.15509926, 17.39302, 3.6827166, 0.76351553, 0.15021779, 15.609284, 3.453064, 0.72047055, 0.14504503, 13.938779, 3.2299175, 0.67823553, 0.13964263, 12.378118, 3.0137942, 0.6369555, 0.13406663, 10.923679, 2.8051126, 0.596754, 0.12836772, 9.571656, 2.6042035, 0.55773467, 0.1225916, 8.318097, 2.4113164, 0.51998276, 0.11677924, 7.1589427, 2.2266283, 0.48356685, 0.11096723, 6.090062, 2.0502505, 0.4485405, 0.10518803, 5.107285, 1.882235, 0.41494337, 0.09947026},
		'{-41.919586, -6.134276, -1.1871881, -0.17252678, -38.91142, -5.896479, -1.150203, -0.17413771, -36.023823, -5.65244, -1.1109434, -0.1745937, -33.25938, -5.404225, -1.0698845, -0.17402205, -30.619717, -5.1536913, -1.0274582, -0.17254148, -28.105562, -4.902501, -0.98405546, -0.17026244, -25.716866, -4.6521325, -0.9400288, -0.16728744, -23.452885, -4.403894, -0.89569455, -0.16371135, -21.31226, -4.158933, -0.8513352, -0.15962176, -19.29309, -3.9182527, -0.80720174, -0.15509926, -17.39302, -3.6827166, -0.76351553, -0.15021779, -15.609284, -3.453064, -0.72047055, -0.14504503, -13.938779, -3.2299175, -0.67823553, -0.13964263, -12.378118, -3.0137942, -0.6369555, -0.13406663, -10.923679, -2.8051126, -0.596754, -0.12836772, -9.571656, -2.6042035, -0.55773467, -0.1225916, -8.318097, -2.4113164, -0.51998276, -0.11677924, -7.1589427, -2.2266283, -0.48356685, -0.11096723, -6.090062, -2.0502505, -0.4485405, -0.10518803, -5.107285, -1.882235, -0.41494337, -0.09947026}};
	localparam real hf[0:1599] = {0.041745532, -0.00026604868, -0.00034630258, 4.1323233e-06, 0.041479833, -0.0007946557, -0.0003372517, 1.2257965e-05, 0.04095213, -0.0013130015, -0.0003194019, 1.9984922e-05, 0.0401692, -0.0018145759, -0.0002931879, 2.7086931e-05, 0.039140992, -0.0022931986, -0.00025920154, 3.337239e-05, 0.037880436, -0.0027431194, -0.00021817042, 3.868457e-05, 0.036403213, -0.003159104, -0.00017093598, 4.2901294e-05, 0.034727477, -0.003536509, -0.000118431104, 4.593421e-05, 0.032873552, -0.0038713403, -6.1657694e-05, 4.7727583e-05, 0.030863572, -0.004160301, -1.6646208e-06, 4.825672e-05, 0.028721146, -0.0044008205, 6.0473703e-05, 4.752605e-05, 0.026470983, -0.004591076, 0.0001236779, 4.556689e-05, 0.024138512, -0.0047299964, 0.000186883, 4.2434967e-05, 0.021749513, -0.0048172553, 0.00024905644, 3.8207734e-05, 0.019329745, -0.004853251, 0.00030921455, 3.2981523e-05, 0.016904594, -0.0048390776, 0.0003664372, 2.6868596e-05, 0.014498732, -0.0047764857, 0.0004198807, 1.999414e-05, 0.012135801, -0.004667831, 0.00046878876, 1.2493248e-05, 0.009838127, -0.0045160227, 0.0005125013, 4.507928e-06, 0.007626455, -0.004324457, 0.00055046135, -3.8158023e-06, 0.0055197245, -0.004096951, 0.00058222, -1.2330718e-05, 0.0035348753, -0.003837672, 0.0006074391, -2.0891037e-05, 0.0016866917, -0.0035510648, 0.00062589237, -2.9354893e-05, -1.2317819e-05, -0.0032417742, 0.00063746434, -3.7586593e-05, -0.001552002, -0.002914573, 0.00064214785, -4.545867e-05, -0.0029246125, -0.002574287, 0.0006400397, -5.2853655e-05, -0.004124812, -0.0022257238, 0.00063133496, -5.966562e-05, -0.0051496476, -0.001873606, 0.0006163203, -6.580144e-05, -0.0059984946, -0.0015225053, 0.0005953654, -7.118177e-05, -0.006672962, -0.0011767856, 0.0005689144, -7.574178e-05, -0.0071767787, -0.0008405481, 0.00053747586, -7.943157e-05, -0.007515648, -0.00051758514, 0.0005016126, -8.221639e-05, -0.0076970835, -0.00021133904, 0.00046193085, -8.407655e-05, -0.0077302256, 7.513145e-05, 0.00041906952, -8.500711e-05, -0.0076256413, 0.00033917773, 0.00037368925, -8.5017375e-05, -0.0073951166, 0.00057858083, 0.00032646157, -8.4130144e-05, -0.0070514353, 0.00079156365, 0.0002780587, -8.238085e-05, -0.006608159, 0.0009767965, 0.00022914326, -7.9816455e-05, -0.0060794014, 0.0011333951, 0.00018035919, -7.649427e-05, -0.0054796096, 0.0012609136, 0.00013232288, -7.248068e-05, -0.0048233466, 0.0013593294, 8.5615306e-05, -6.784975e-05, -0.004125083, 0.0014290254, 4.0775074e-05, -6.26818e-05, -0.0033990038, 0.0014707638, -1.707661e-06, -5.7061898e-05, -0.0026588228, 0.0014856587, -4.1396266e-05, -5.1078445e-05, -0.0019176156, 0.0014751424, -7.791166e-05, -4.482169e-05, -0.0011876696, 0.0014409306, -0.00011093531, -3.8382303e-05, -0.00048035113, 0.0013849838, -0.0001402112, -3.1850017e-05, 0.00019400618, 0.0013094669, -0.0001655468, -2.5312353e-05, 0.0008261942, 0.0012167093, -0.00018681296, -1.8853398e-05, 0.0014082015, 0.0011091623, -0.0002039431, -1.2552735e-05, 0.0019332647, 0.0009893584, -0.00021693118, -6.4844567e-06, 0.0023958979, 0.00085987063, -0.00022582914, -7.1631774e-07, 0.0027919041, 0.0007232735, -0.00023074354, 4.690981e-06, 0.0031183658, 0.0005821055, -0.00023183145, 9.6843705e-06, 0.0033736182, 0.00043883413, -0.0002292959, 1.42188555e-05, 0.0035572064, 0.000295824, -0.00022338083, 1.8257813e-05, 0.003669825, 0.00015530705, -0.00021436562, 2.1773152e-05, 0.0037132464, 1.9357152e-05, -0.00020255946, 2.4745343e-05, 0.0036902358, -0.00011013236, -0.00018829544, 2.7163322e-05, 0.0036044552, -0.0002314672, -0.00017192465, 2.9024262e-05, 0.0034603616, -0.00034316684, -0.0001538102, 3.0333247e-05, 0.003263096, -0.0004439754, -0.00013432144, 3.1102838e-05, 0.00301837, -0.0005328687, -0.00011382835, 3.135254e-05, 0.0027323477, -0.0006090576, -9.269606e-05, 3.1108226e-05, 0.0024115301, -0.0006719875, -7.127988e-05, 3.040143e-05, 0.0020626367, -0.00072133465, -4.9920596e-05, 2.9268664e-05, 0.0016924929, -0.0007569995, -2.8940236e-05, 2.7750637e-05, 0.0013079197, -0.00077909604, -8.6383125e-06, 2.5891475e-05, 0.0009156302, -0.0007879401, 1.0711427e-05, 2.3737924e-05, 0.0005221323, -0.00078403373, 2.8863718e-05, 2.133855e-05, 0.00013363991, -0.00076804834, 4.5603938e-05, 1.8742943e-05, -0.00024400756, -0.0007408064, 6.0749724e-05, 1.6000959e-05, -0.0006054154, -0.0007032612, 7.4152034e-05, 1.3161975e-05, -0.00094569376, -0.0006564759, 8.569567e-05, 1.027421e-05, -0.0012605077, -0.00060160225, 9.529925e-05, 7.3840665e-06, -0.0015461156, -0.00053985894, 0.00010291475, 4.5355578e-06, -0.0017993973, -0.00047250945, 0.00010852651, 1.7697766e-06, -0.0020178712, -0.00040084135, 0.00011214983, -8.7555475e-07, -0.0021997013, -0.0003261454, 0.000113829214, -3.3664708e-06, -0.0023436933, -0.0002496961, 0.00011363622, -5.6730714e-06, -0.002449283, -0.00017273327, 0.00011166705, -7.769757e-06, -0.0025165125, -9.644509e-05, 0.00010803987, -9.6353915e-06, -0.0025460033, -2.1952763e-05, 0.00010289197, -1.1253385e-05, -0.002538917, 4.970307e-05, 9.637675e-05, -1.26117175e-05, -0.002496913, 0.00011757407, 8.8660614e-05, -1.3702878e-05, -0.0024220997, 0.00018081395, 7.9919846e-05, -1.4523757e-05, -0.0023169818, 0.00023868626, 7.0337504e-05, -1.50754695e-05, -0.002184403, 0.00029057014, 6.0100305e-05, -1.536312e-05, -0.0020274878, 0.00033596397, 4.9395687e-05, -1.5395543e-05, -0.0018495816, 0.00037448722, 3.8408944e-05, -1.518496e-05, -0.0016541894, 0.00040588036, 2.7320575e-05, -1.4746654e-05, -0.0014449162, 0.00043000278, 1.6303806e-05, -1.4098571e-05, -0.0012254084, 0.00044682936, 5.5223563e-06, -1.3260929e-05, -0.0009992969, 0.00045644512, -4.871546e-06, -1.2255797e-05, -0.0007701439, 0.00045903886, -1.4738881e-05, -1.1106677e-05, -0.00054139306, 0.0004548951, -2.3955274e-05, -9.838082e-06, -0.00031632345, 0.0004443856, -3.2412143e-05, -8.475117e-06, -9.800861e-05, 0.00042795928, -4.0017552e-05, -7.043077e-06, 0.00011071963, 0.00040613202, -4.669678e-05, -5.5670557e-06, 0.00030730182, 0.00037947576, -5.23926e-05, -4.0715845e-06, 0.00048947614, 0.00034860722, -5.706529e-05, -2.5802892e-06, 0.00065529795, 0.00031417652, -6.069237e-05, -1.1155827e-06, 0.0008031538, 0.0002768561, -6.326812e-05, 3.016111e-07, 0.00093176943, 0.00023732937, -6.480283e-05, 1.652098e-06, 0.001040213, 0.00019628023, -6.532189e-05, 2.9186162e-06, 0.0011278928, 0.00015438274, -6.486468e-05, 4.086e-06, 0.0011945489, 0.000112291564, -6.34833e-05, 5.141305e-06, 0.001240243, 7.0633265e-05, -6.124117e-05, 6.073893e-06, 0.0012653406, 2.9998188e-05, -5.821157e-05, 6.87548e-06, 0.0012704922, -9.066478e-06, -5.4476033e-05, 7.5401445e-06, 0.0012566097, -4.6062818e-05, -5.012275e-05, 8.064302e-06, 0.0012248404, -8.0547215e-05, -4.5244935e-05, 8.446648e-06, 0.0011765393, -0.00011213436, -3.9939183e-05, 8.688061e-06, 0.0011132385, -0.00014050014, -3.4303874e-05, 8.791489e-06, 0.0010366167, -0.00016538358, -2.8437618e-05, 8.761804e-06, 0.0009484669, -0.00018658763, -2.2437784e-05, 8.605636e-06, 0.00085066474, -0.00020397906, -1.639909e-05, 8.33119e-06, 0.00074513664, -0.00021748741, -1.0412333e-05, 7.948044e-06, 0.00063382904, -0.00022710294, -4.563222e-06, 7.4669465e-06, 0.0005186786, -0.00023287392, 1.0686539e-06, 6.8995923e-06, 0.000401584, -0.00023490313, 6.410718e-06, 6.2584086e-06, 0.00028437976, -0.0002333437, 1.1398149e-05, 5.55633e-06, 0.00016881226, -0.0002283944, 1.597447e-05, 4.8065845e-06, 5.6518104e-05, -0.00022029456, 2.0091995e-05, 4.0224795e-06, -5.0994746e-05, -0.00020931849, 2.3712108e-05, 3.2172018e-06, -0.00015236306, -0.0001957698, 2.680541e-05, 2.4036246e-06, -0.00024638147, -0.00017997542, 2.9351706e-05, 1.5941337e-06, -0.00033201274, -0.00016227973, 3.1339867e-05, 8.004638e-07, -0.00040839482, -0.00014303849, 3.2767566e-05, 3.3556752e-08, -0.00047484526, -0.00012261311, 3.3640874e-05, -6.9656414e-07, -0.0005308625, -0.00010136495, 3.397379e-05, -1.380899e-06, -0.0005761245, -7.965005e-05, 3.3787623e-05, -2.0115558e-06, -0.00061048503, -5.7814017e-05, 3.3110355e-05, -2.581815e-06, -0.0006339667, -3.6187455e-05, 3.197588e-05, -3.0861731e-06, -0.0006467532, -1.5081782e-05, 3.0423233e-05, -3.5203661e-06, -0.00064917805, 5.2144746e-06, 2.8495751e-05, -3.8813732e-06, -0.0006417128, 2.443884e-05, 2.624024e-05, -4.167402e-06, -0.00062495307, 4.2357522e-05, 2.3706087e-05, -4.3778564e-06, -0.0005996038, 5.8767506e-05, 2.0944432e-05, -4.5132883e-06, -0.0005664634, 7.349806e-05, 1.8007306e-05, -4.5753336e-06, -0.00052640727, 8.641171e-05, 1.4946819e-05, -4.5666357e-06, -0.00048037132, 9.7404685e-05, 1.1814389e-05, -4.490758e-06, -0.00042933473, 0.00010640679, 8.6600085e-06, -4.3520886e-06, -0.00037430358, 0.000113380855, 5.5315704e-06, -4.155732e-06, -0.0003162945, 0.00011832167, 2.4742617e-06, -3.907401e-06, -0.00025631895, 0.000121254496, -4.6997877e-07, -3.613304e-06, -0.00019536859, 0.00012223326, -3.2629237e-06, -3.2800256e-06, -0.00013440137, 0.00012133831, -5.870446e-06, -2.914413e-06, -7.432899e-05, 0.000118673976, -8.262828e-06, -2.5234622e-06, -1.600553e-05, 0.00011436584, -1.0414987e-05, -2.1142048e-06, 3.9782444e-05, 0.00010855784, -1.2306627e-05, -1.6936041e-06, 9.232428e-05, 0.00010140926, -1.3922302e-05, -1.2684541e-06, 0.00014099214, 9.309159e-05, -1.5251419e-05, -8.45287e-07, 0.00018524638, 8.378541e-05, -1.6288155e-05, -4.302888e-07, 0.00022463918, 7.3677234e-05, -1.7031312e-05, -2.9224458e-08, 0.0002588169, 6.29565e-05, -1.7484113e-05, 3.5262744e-07, 0.0002875207, 5.1812534e-05, -1.7653942e-05, 7.105295e-07, 0.0003105858, 4.043184e-05, -1.7552025e-05, 1.0403297e-06, 0.00032793934, 2.8995384e-05, -1.7193088e-05, 1.3384947e-06, 0.0003395971, 1.7676197e-05, -1.659496e-05, 1.6021322e-06, 0.000345659, 6.6371917e-06, -1.5778161e-05, 1.8290033e-06, 0.0003463033, -3.970771e-06, -1.4765471e-05, 2.0175235e-06, 0.0003417805, -1.40105485e-05, -1.3581472e-05, 2.166755e-06, 0.00033240582, -2.3360086e-05, -1.2252103e-05, 2.2763893e-06, 0.00031855155, -3.1913507e-05, -1.08042095e-05, 2.3467212e-06, 0.0003006387, -3.9581897e-05, -9.265097e-06, 2.378615e-06, 0.00027912838, -4.6293808e-05, -7.662104e-06, 2.3734647e-06, 0.00025451303, -5.1995485e-05, -6.022192e-06, 2.333147e-06, 0.00022730745, -5.6650795e-05, -4.3715686e-06, 2.2599704e-06, 0.0001980403, -6.0240916e-05, -2.7353294e-06, 2.15662e-06, 0.00016724532, -6.276379e-05, -1.1371408e-06, 2.0260989e-06, 0.0001354533, -6.4233325e-05, 4.010435e-07, 1.8716687e-06, 0.00010318427, -6.467843e-05, 1.8592249e-06, 1.6967887e-06, 7.094028e-05, -6.414185e-05, 3.2195635e-06, 1.5050541e-06, 3.9198825e-05, -6.267888e-05, 4.466538e-06, 1.3001369e-06, 8.406919e-06, -6.035591e-05, 5.587065e-06, 1.0857268e-06, -2.1024085e-05, -5.7248908e-05, 6.570575e-06, 8.65476e-07, -4.872289e-05, -5.3441847e-05, 7.409048e-06, 6.4294665e-07, -7.436183e-05, -4.9025046e-05, 8.097009e-06, 4.2156222e-07, -9.765966e-05, -4.4093536e-05, 8.631489e-06, 2.0456325e-07, -0.00011838346, -3.874541e-05, 9.011942e-06, -5.031821e-09, -0.0001363498, -3.3080214e-05, 9.240142e-06, -2.0446087e-07, -0.00015142508, -2.7197406e-05, 9.320041e-06, -3.9124672e-07, -0.00016352505, -2.1194879e-05, 9.257604e-06, -5.6322017e-07, -0.00017261377, -1.51675795e-05, 9.060629e-06, -7.185373e-07, -0.00017870174, -9.2062355e-06, 8.738533e-06, -8.5569127e-07, -0.00018184353, -3.3962156e-06, 8.302143e-06, -9.735182e-07, -0.00018213484, 2.1834817e-06, 7.7634595e-06, -1.0711982e-06, -0.00017970912, 7.4610953e-06, 7.135425e-06, -1.1482504e-06, -0.00017473368, 1.237282e-05, 6.4316873e-06, -1.2045243e-06, -0.00016740568, 1.6863367e-05, 5.666358e-06, -1.2401855e-06, -0.00015794765, 2.0886377e-05, 4.853784e-06, -1.2556984e-06, -0.00014660307, 2.440468e-05, 4.0083223e-06, -1.2518045e-06, -0.00013363162, 2.7390399e-05, 3.1441236e-06, -1.229498e-06, -0.00011930462, 2.9824914e-05, 2.2749355e-06, -1.1899991e-06, -0.00010390044, 3.1698703e-05, 1.4139143e-06, -1.1347245e-06, -8.769998e-05, 3.301103e-05, 5.734608e-07, -1.065257e-06, -7.0982365e-05, 3.376954e-05, -2.3493e-07, -9.833144e-07, -5.4020962e-05, 3.398973e-05, -1.0007943e-06, -8.9071654e-07, -3.7079502e-05, 3.3694363e-05, -1.714806e-06, -7.893539e-07, -2.0408694e-05, 3.2912747e-05, -2.3688601e-06, -6.811561e-07, -4.24309e-06, 3.168001e-05, -2.9561345e-06, -5.6806107e-07, 1.1201599e-05, 3.003628e-05, -3.4711288e-06, -4.519859e-07, 2.5730804e-05, 2.8025852e-05, -3.9096826e-06, -3.3479944e-07, 3.917297e-05, 2.569633e-05, -4.268973e-06, -2.1829676e-07, 5.1380986e-05, 2.3097758e-05, -4.547491e-06, -1.041761e-07, 6.223319e-05, 2.0281763e-05, -4.7450003e-06, 5.981753e-09, 7.163397e-05, 1.7300701e-05, -4.862482e-06, 1.107313e-07, 7.9513884e-05, 1.4206852e-05, -4.902057e-06, 2.0877722e-07, 8.5829444e-05, 1.1051647e-05, -4.8669017e-06, 2.9898644e-07, 9.0562535e-05, 7.884938e-06, -4.761151e-06, 3.8039704e-07, 9.371941e-05, 4.754341e-06, -4.589788e-06, 4.5222438e-07, 9.532947e-05, 1.7046308e-06, -4.35853e-06, 5.1386417e-07, 9.5443655e-05, -1.2227831e-06, -4.073709e-06, 5.648927e-07, 9.413267e-05, -3.990312e-06, -3.7421453e-06, 6.050644e-07, 9.148501e-05, -6.5645604e-06, -3.3710255e-06, 6.3430696e-07, 8.760472e-05, -8.916621e-06, -2.9677767e-06, 6.52714e-07, 8.260916e-05, -1.1022283e-05, -2.539944e-06, 6.605356e-07, 7.662656e-05, -1.2862173e-05, -2.0950731e-06, 6.581671e-07, 6.9793634e-05, -1.4421801e-05, -1.6405986e-06, 6.461362e-07, 6.2253115e-05, -1.5691545e-05, -1.183738e-06, 6.250886e-07, 5.4151365e-05, -1.6666554e-05, -7.313957e-07, 5.957729e-07, 4.563598e-05, -1.7346594e-05, -2.900748e-07, 5.590244e-07, 3.6853584e-05, -1.7735827e-05, 1.3419942e-07, 5.157483e-07, 2.794767e-05, -1.7842533e-05, 5.359465e-07, 4.6690323e-07, 1.9056624e-05, -1.767879e-05, 9.102856e-07, 4.1348426e-07, 1.0311924e-05, -1.726012e-05, 1.2529792e-06, 3.5650626e-07, 1.836507e-06, -1.660507e-05, 1.5604652e-06, 2.9698796e-07, -6.2566364e-06, -1.5734817e-05, 1.8298765e-06, 2.3593658e-07, -1.3865663e-05, -1.4672701e-05, 2.0590508e-06, 1.7433346e-07, -2.0900854e-05, -1.3443791e-05, 2.246528e-06, 1.13120706e-07, -2.7285358e-05, -1.20744235e-05, 2.391539e-06, 5.318905e-08, -3.295571e-05, -1.0591746e-05, 2.4939823e-06, -4.6328443e-09, -3.786214e-05, -9.02328e-06, 2.5543943e-06, -5.9587748e-08, -4.1968633e-05, -7.396488e-06, 2.5739098e-06, -1.1099764e-07, -4.5252804e-05, -5.738375e-06, 2.554217e-06, -1.5826997e-07, -4.7705584e-05, -4.0751033e-06, 2.497505e-06, -2.009023e-07, -4.9330694e-05, -2.4316482e-06, 2.406407e-06, -2.3848548e-07, -5.0143983e-05, -8.314821e-07, 2.2839404e-06, -2.7070516e-07, -5.01726e-05, 7.037013e-07, 2.1334424e-06, -2.973419e-07, -4.9454047e-05, 2.1542228e-06, 1.9585061e-06, -3.1826983e-07, -4.8035115e-05, 3.502613e-06, 1.7629134e-06, -3.3345404e-07, -4.597075e-05, 4.733766e-06, 1.5505706e-06, -3.4294666e-07, -4.3322838e-05, 5.835049e-06, 1.3254444e-06, -3.4688188e-07, -4.015894e-05, 6.7963683e-06, 1.091499e-06, -3.4546997e-07, -3.655102e-05, 7.6102024e-06, 8.526388e-07, -3.3899056e-07, -3.2574175e-05, 8.271582e-06, 6.126518e-07, -3.2778505e-07, -2.8305343e-05, 8.778047e-06, 3.751598e-07, -3.1224855e-07, -2.3822091e-05, 9.129557e-06, 1.435725e-07, -2.9282148e-07, -1.9201418e-05, 9.328378e-06, -7.8953136e-08, -2.6998077e-07, -1.4518649e-05, 9.378936e-06, -2.895475e-07, -2.44231e-07, -9.846386e-06, 9.287646e-06, -4.856571e-07, -2.160956e-07, -5.2535684e-06, 9.062723e-06, -6.650671e-07, -1.8610817e-07, -8.0462104e-07, 8.713968e-06, -8.259181e-07, -1.5480401e-07, 3.4412838e-06, 8.252551e-06, -9.667165e-07, -1.2271214e-07, 7.4308523e-06, 7.690779e-06, -1.0863387e-06, -9.034764e-08, 1.1117177e-05, 7.04185e-06, -1.1840305e-06, -5.820481e-08, 1.4460125e-05, 6.3196244e-06, -1.2593999e-06, -2.6750717e-08, 1.7426608e-05, 5.5383794e-06, -1.312406e-06, 3.5803926e-09, 1.999073e-05, 4.71258e-06, -1.3433419e-06, 3.2391956e-08, 2.213383e-05, 3.8566545e-06, -1.3528147e-06, 5.932917e-08, 2.3844408e-05, 2.984781e-06, -1.3417213e-06, 8.408225e-08, 2.5117946e-05, 2.1106891e-06, -1.3112208e-06, 1.0638886e-07, 2.595664e-05, 1.2474783e-06, -1.2627047e-06, 1.2603569e-07, 2.6369045e-05, 4.0745232e-07, -1.1977652e-06, 1.4285932e-07, 2.6369638e-05, -3.980239e-07, -1.1181614e-06, 1.5674614e-07, 2.5978317e-05, -1.1586486e-06, -1.0257855e-06, 1.6763174e-07, 2.521984e-05, -1.8652848e-06, -9.2262803e-07, 1.754994e-07, 2.4123232e-05, -2.5100396e-06, -8.1074336e-07, 1.8037807e-07, 2.2721133e-05, -3.0863212e-06, -6.9221653e-07, 1.8233975e-07, 2.104915e-05, -3.5888745e-06, -5.691303e-07, 1.8149628e-07, 1.9145182e-05, -4.0137943e-06, -4.4353462e-07, 1.7799583e-07, 1.7048738e-05, -4.358518e-06, -3.174176e-07, 1.7201887e-07, 1.4800284e-05, -4.6217983e-06, -1.92679e-07, 1.6377396e-07, 1.2440583e-05, -4.80366e-06, -7.1106214e-08, 1.5349329e-07, 1.0010085e-05, -4.9053356e-06, 4.564679e-08, 1.414281e-07, 7.5483367e-06, -4.9291907e-06, 1.5607766e-07, 1.2784398e-07, 5.0934354e-06, -4.8786324e-06, 2.5885066e-07, 1.1301628e-07, 2.6815364e-06, -4.75801e-06, 3.5280843e-07, 9.7225495e-08, 3.4640763e-07, -4.5725033e-06, 4.3698057e-07, 8.075291e-08, -1.8809568e-06, -4.328006e-06, 5.1058913e-07, 6.3876314e-08, -3.9726624e-06, -4.031004e-06, 5.730506e-07, 4.68661e-08, -5.9041804e-06, -3.6884505e-06, 6.239756e-07, 2.9981543e-08, -7.654547e-06, -3.3076383e-06, 6.631648e-07, 1.3467543e-08, -9.206506e-06, -2.8960771e-06, 6.906032e-07, -2.448364e-09, -1.0546583e-05, -2.4613707e-06, 7.06451e-07, -1.7558524e-08, -1.1665106e-05, -2.011099e-06, 7.1103284e-07, -3.16773e-08, -1.2556163e-05, -1.5527066e-06, 7.048254e-07, -4.4642764e-08, -1.32175055e-05, -1.0933995e-06, 6.884425e-07, -5.6317965e-08, -1.3650413e-05, -6.400486e-07, 6.626196e-07, -6.659174e-08, -1.3859495e-05, -1.9910387e-07, 6.2819674e-07, -7.5379134e-08, -1.3852466e-05, 2.2348063e-07, 5.861014e-07, -8.26214e-08, -1.36398785e-05, 6.223117e-07, 5.3733015e-07, -8.828558e-08, -1.3234832e-05, 9.926099e-07, 4.8293055e-07, -9.236379e-08, -1.2652653e-05, 1.3302508e-06, 4.2398335e-07, -9.487207e-08, -1.1910556e-05, 1.6317953e-06, 3.6158445e-07, -9.584904e-08, -1.1027305e-05, 1.8945062e-06, 2.968282e-07, -9.535421e-08, -1.0022853e-05, 2.1163567e-06, 2.3079103e-07, -9.3466085e-08, -8.917988e-06, 2.2960246e-06, 1.6451636e-07, -9.028008e-08, -7.733988e-06, 2.432879e-06, 9.9000744e-08, -8.59063e-08, -6.4922774e-06, 2.5269558e-06, 3.5181213e-08, -8.046717e-08, -5.214102e-06, 2.5789248e-06, -2.607566e-08, -7.4095034e-08, -3.920223e-06, 2.5900495e-06, -8.398331e-08, -6.6929715e-08, -2.6306316e-06, 2.5621393e-06, -1.3784297e-07, -5.9116044e-08, -1.3642878e-06, 2.497496e-06, -1.8704985e-07, -5.080151e-08, -1.3889007e-07, 2.3988569e-06, -2.3109749e-07, -4.2133905e-08, 1.0293274e-06, 2.2693312e-06, -2.6958065e-07, -3.325912e-08, 2.1257656e-06, 2.1123374e-06, -3.021964e-07, -2.4319084e-08, 3.1375978e-06, 1.9315373e-06, -3.2874362e-07, -1.5449821e-08, 4.0538753e-06, 1.7307689e-06, -3.491211e-07, -6.779738e-09, 4.8655984e-06, 1.5139818e-06, -3.6332432e-07, 1.5719323e-09, 5.565757e-06, 1.2851727e-06, -3.7144062e-07, 9.496452e-09, 6.149339e-06, 1.0483236e-06, -3.7364367e-07, 1.689669e-08, 6.6133052e-06, 8.0734367e-07, -3.7018663e-07, 2.3688003e-08, 6.956543e-06, 5.660143e-07, -3.6139448e-07, 2.9798889e-08, 7.1797876e-06, 3.2793946e-07, -3.476559e-07, 3.5171418e-08, 7.285522e-06, 9.650032e-08, -3.294142e-07, 3.976144e-08, 7.2778557e-06, -1.2518392e-07, -3.0715825e-07, 4.3538552e-08, 7.162385e-06, -3.342899e-07, -2.814129e-07, 4.648593e-08, 6.9460384e-06, -5.283177e-07, -2.527295e-07, 4.859987e-08, 6.636909e-06, -7.051124e-07, -2.2167647e-07, 4.9889252e-08, 6.244076e-06, -8.628794e-07, -1.8882989e-07, 5.0374776e-08, 5.7774255e-06, -1.0001936e-06, -1.5476468e-07, 5.0088094e-08, 5.247463e-06, -1.116003e-06, -1.200461e-07, 4.907079e-08, 4.6651253e-06, -1.2096259e-06, -8.522175e-08, 4.7373316e-08, 4.041601e-06, -1.2807433e-06, -5.081436e-08, 4.5053785e-08, 3.3881486e-06, -1.3293862e-06, -1.7315188e-08, 4.2176744e-08, 2.7159272e-06, -1.3559182e-06, 1.4821778e-08, 3.8811912e-08, 2.0358364e-06, -1.361014e-06, 4.5184727e-08, 3.5032883e-08, 1.3583644e-06, -1.3456342e-06, 7.340813e-08, 3.0915857e-08, 6.9345475e-07, -1.3109972e-06, 9.917594e-08, 2.6538357e-08, 5.038252e-08, -1.2585489e-06, 1.2222388e-07, 2.197805e-08, -5.6234967e-07, -1.1899299e-06, 1.4234087e-07, 1.731155e-08, -1.1371013e-06, -1.106942e-06, 1.5936959e-07, 1.2613351e-08, -1.6671659e-06, -1.0115133e-06, 1.7320627e-07, 7.954819e-09, -2.1468254e-06, -9.0566357e-07, 1.8379957e-07, 3.4032754e-09, -2.571387e-06, -7.9147003e-07, 1.9114884e-07, -9.788003e-10, -2.9372043e-06, -6.710333e-07, 1.9530167e-07, -5.134469e-09, -3.2416801e-06, -5.464454e-07, 1.9635088e-07, -9.0129095e-09, -3.4832542e-06, -4.1975866e-07, 1.9443092e-07, -1.2569879e-08, -3.6613771e-06, -2.9295762e-07, 1.8971389e-07, -1.576805e-08, -3.776469e-06, -1.6793253e-07, 1.8240512e-07, -1.8577236e-08, -3.8298663e-06, -4.6455742e-08, 1.7273852e-07, -2.0974484e-08, -3.823758e-06, 6.983869e-08, 1.609718e-07, -2.2944084e-08, -3.7611119e-06, 1.794728e-07, 1.4738134e-07, -2.4477433e-08, -3.6455922e-06, 2.8113908e-07, 1.3225736e-07, -2.5572833e-08, -3.4814725e-06, 3.737116e-07, 1.1589875e-07, -2.6235176e-08, -3.273541e-06, 4.562541e-07, 9.860837e-08, -2.6475552e-08, -3.0270073e-06, 5.280246e-07, 8.068825e-08, -2.6310792e-08, -2.7474011e-06, 5.884772e-07, 6.243519e-08, -2.5762928e-08, -2.4404778e-06, 6.372605e-07, 4.4136584e-08, -2.4858627e-08, -2.1121195e-06, 6.7421354e-07, 2.6066619e-08, -2.3628562e-08, -1.768243e-06, 6.993591e-07, 8.482815e-09, -2.2106766e-08, -1.4147099e-06, 7.1289423e-07, -8.376974e-09, -2.032996e-08, -1.0572415e-06, 7.1517906e-07, -2.429716e-08, -1.8336882e-08, -7.013413e-07, 7.0672354e-07, -3.908654e-08, -1.6167615e-08, -3.522233e-07, 6.881726e-07, -5.2579967e-08, -1.3862916e-08, -1.4748624e-08, 6.6029e-07, -6.4639536e-08, -1.146359e-08, 3.066297e-07, 6.239414e-07, -7.515533e-08, -9.009873e-09, 6.079131e-07, 5.800763e-07, -8.4045666e-08, -6.5408656e-09, 8.85595e-07, 5.2971006e-07, -9.125701e-08, -4.0940042e-09, 1.1366892e-06, 4.7390563e-07, -9.676333e-08, -1.7045872e-09, 1.3587492e-06, 4.1375532e-07, -1.0056523e-07, 5.946482e-10, 1.5498778e-06, 3.5036328e-07, -1.02688595e-07, 2.7738878e-09, 1.7087299e-06, 2.8482845e-07, -1.0318301e-07, 4.806542e-09, 1.8345047e-06, 2.1822848e-07, -1.021199e-07, 6.669485e-09, 1.926932e-06, 1.5160478e-07, -9.959034e-08, 8.343233e-09, 1.9862505e-06, 8.594872e-08, -9.570284e-08, 9.812055e-09, 2.0131788e-06, 2.2189392e-08, -9.058082e-08, 1.1064026e-08, 2.0088828e-06, -3.881723e-08, -8.43601e-08, 1.2091022e-08, 1.9749357e-06, -9.629747e-08, -7.718627e-08, 1.2888656e-08, 1.913276e-06, -1.4956747e-07, -6.921202e-08, 1.345616e-08, 1.8261597e-06, -1.98039e-07, -6.059457e-08, 1.3796225e-08, 1.7161124e-06, -2.4122363e-07, -5.149311e-08, 1.3914792e-08, 1.5858784e-06, -2.7873506e-07, -4.206631e-08, 1.3820808e-08, 1.4383693e-06, -3.1029006e-07, -3.2470016e-08, 1.3525944e-08, 1.2766128e-06, -3.3570754e-07, -2.2855051e-08, 1.3044296e-08, 1.103702e-06, -3.549065e-07, -1.336523e-08, 1.2392054e-08, 9.2274604e-07, -3.6790215e-07, -4.135552e-09, 1.1587158e-08, 7.3682355e-07, -3.748013e-07, 4.709376e-09, 1.0648952e-08, 5.489381e-07, -3.757961e-07, 1.3056691e-08, 9.5978265e-09, 3.619772e-07, -3.7115723e-07, 2.080638e-08, 8.454863e-09, 1.7867491e-07, -3.6122603e-07, 2.7872154e-08, 7.24149e-09, 1.5789132e-09, -3.4640595e-07, 3.418205e-08, 5.979147e-09, -1.6697864e-07, -3.2715363e-07, 3.9678834e-08, 4.688963e-09, -3.2490524e-07, -3.039695e-07, 4.4320114e-08, 3.391461e-09, -4.7036752e-07, -2.7738824e-07, 4.8078263e-08, 2.1062794e-09, -6.0180605e-07, -2.4796915e-07, 5.0940116e-08, 8.5192514e-10, -7.1794517e-07, -2.1628675e-07, 5.2906476e-08, -3.5444864e-10, -8.1779837e-07, -1.8292133e-07, 5.3991403e-08, -1.4972308e-09, -9.0066885e-07, -1.4845017e-07, 5.4221392e-08, -2.5625104e-09, -9.66146e-07, -1.134391e-07, 5.363435e-08, -3.5382006e-09, -1.0140974e-06, -7.8434596e-08, 5.227851e-08, -4.414131e-09, -1.0446577e-06, -4.3956618e-08, 5.0211185e-08, -5.182105e-09, -1.0582135e-06, -1.0492179e-08, 4.7497505e-08, -5.8359273e-09, -1.0553852e-06, 2.1510338e-08, 4.420905e-08, -6.371399e-09, -1.0370072e-06, 5.1645944e-08, 4.0422485e-08, -6.7862826e-09, -1.0041043e-06, 7.955698e-08, 3.621818e-08, -7.080242e-09, -9.578679e-07, 1.04936156e-07, 3.167881e-08, -7.254754e-09, -8.9962964e-07, 1.2752865e-07, 2.688805e-08, -7.3129995e-09};
	localparam real hb[0:1599] = {0.041745532, 0.00026604868, -0.00034630258, -4.1323233e-06, 0.041479833, 0.0007946557, -0.0003372517, -1.2257965e-05, 0.04095213, 0.0013130015, -0.0003194019, -1.9984922e-05, 0.0401692, 0.0018145759, -0.0002931879, -2.7086931e-05, 0.039140992, 0.0022931986, -0.00025920154, -3.337239e-05, 0.037880436, 0.0027431194, -0.00021817042, -3.868457e-05, 0.036403213, 0.003159104, -0.00017093598, -4.2901294e-05, 0.034727477, 0.003536509, -0.000118431104, -4.593421e-05, 0.032873552, 0.0038713403, -6.1657694e-05, -4.7727583e-05, 0.030863572, 0.004160301, -1.6646208e-06, -4.825672e-05, 0.028721146, 0.0044008205, 6.0473703e-05, -4.752605e-05, 0.026470983, 0.004591076, 0.0001236779, -4.556689e-05, 0.024138512, 0.0047299964, 0.000186883, -4.2434967e-05, 0.021749513, 0.0048172553, 0.00024905644, -3.8207734e-05, 0.019329745, 0.004853251, 0.00030921455, -3.2981523e-05, 0.016904594, 0.0048390776, 0.0003664372, -2.6868596e-05, 0.014498732, 0.0047764857, 0.0004198807, -1.999414e-05, 0.012135801, 0.004667831, 0.00046878876, -1.2493248e-05, 0.009838127, 0.0045160227, 0.0005125013, -4.507928e-06, 0.007626455, 0.004324457, 0.00055046135, 3.8158023e-06, 0.0055197245, 0.004096951, 0.00058222, 1.2330718e-05, 0.0035348753, 0.003837672, 0.0006074391, 2.0891037e-05, 0.0016866917, 0.0035510648, 0.00062589237, 2.9354893e-05, -1.2317819e-05, 0.0032417742, 0.00063746434, 3.7586593e-05, -0.001552002, 0.002914573, 0.00064214785, 4.545867e-05, -0.0029246125, 0.002574287, 0.0006400397, 5.2853655e-05, -0.004124812, 0.0022257238, 0.00063133496, 5.966562e-05, -0.0051496476, 0.001873606, 0.0006163203, 6.580144e-05, -0.0059984946, 0.0015225053, 0.0005953654, 7.118177e-05, -0.006672962, 0.0011767856, 0.0005689144, 7.574178e-05, -0.0071767787, 0.0008405481, 0.00053747586, 7.943157e-05, -0.007515648, 0.00051758514, 0.0005016126, 8.221639e-05, -0.0076970835, 0.00021133904, 0.00046193085, 8.407655e-05, -0.0077302256, -7.513145e-05, 0.00041906952, 8.500711e-05, -0.0076256413, -0.00033917773, 0.00037368925, 8.5017375e-05, -0.0073951166, -0.00057858083, 0.00032646157, 8.4130144e-05, -0.0070514353, -0.00079156365, 0.0002780587, 8.238085e-05, -0.006608159, -0.0009767965, 0.00022914326, 7.9816455e-05, -0.0060794014, -0.0011333951, 0.00018035919, 7.649427e-05, -0.0054796096, -0.0012609136, 0.00013232288, 7.248068e-05, -0.0048233466, -0.0013593294, 8.5615306e-05, 6.784975e-05, -0.004125083, -0.0014290254, 4.0775074e-05, 6.26818e-05, -0.0033990038, -0.0014707638, -1.707661e-06, 5.7061898e-05, -0.0026588228, -0.0014856587, -4.1396266e-05, 5.1078445e-05, -0.0019176156, -0.0014751424, -7.791166e-05, 4.482169e-05, -0.0011876696, -0.0014409306, -0.00011093531, 3.8382303e-05, -0.00048035113, -0.0013849838, -0.0001402112, 3.1850017e-05, 0.00019400618, -0.0013094669, -0.0001655468, 2.5312353e-05, 0.0008261942, -0.0012167093, -0.00018681296, 1.8853398e-05, 0.0014082015, -0.0011091623, -0.0002039431, 1.2552735e-05, 0.0019332647, -0.0009893584, -0.00021693118, 6.4844567e-06, 0.0023958979, -0.00085987063, -0.00022582914, 7.1631774e-07, 0.0027919041, -0.0007232735, -0.00023074354, -4.690981e-06, 0.0031183658, -0.0005821055, -0.00023183145, -9.6843705e-06, 0.0033736182, -0.00043883413, -0.0002292959, -1.42188555e-05, 0.0035572064, -0.000295824, -0.00022338083, -1.8257813e-05, 0.003669825, -0.00015530705, -0.00021436562, -2.1773152e-05, 0.0037132464, -1.9357152e-05, -0.00020255946, -2.4745343e-05, 0.0036902358, 0.00011013236, -0.00018829544, -2.7163322e-05, 0.0036044552, 0.0002314672, -0.00017192465, -2.9024262e-05, 0.0034603616, 0.00034316684, -0.0001538102, -3.0333247e-05, 0.003263096, 0.0004439754, -0.00013432144, -3.1102838e-05, 0.00301837, 0.0005328687, -0.00011382835, -3.135254e-05, 0.0027323477, 0.0006090576, -9.269606e-05, -3.1108226e-05, 0.0024115301, 0.0006719875, -7.127988e-05, -3.040143e-05, 0.0020626367, 0.00072133465, -4.9920596e-05, -2.9268664e-05, 0.0016924929, 0.0007569995, -2.8940236e-05, -2.7750637e-05, 0.0013079197, 0.00077909604, -8.6383125e-06, -2.5891475e-05, 0.0009156302, 0.0007879401, 1.0711427e-05, -2.3737924e-05, 0.0005221323, 0.00078403373, 2.8863718e-05, -2.133855e-05, 0.00013363991, 0.00076804834, 4.5603938e-05, -1.8742943e-05, -0.00024400756, 0.0007408064, 6.0749724e-05, -1.6000959e-05, -0.0006054154, 0.0007032612, 7.4152034e-05, -1.3161975e-05, -0.00094569376, 0.0006564759, 8.569567e-05, -1.027421e-05, -0.0012605077, 0.00060160225, 9.529925e-05, -7.3840665e-06, -0.0015461156, 0.00053985894, 0.00010291475, -4.5355578e-06, -0.0017993973, 0.00047250945, 0.00010852651, -1.7697766e-06, -0.0020178712, 0.00040084135, 0.00011214983, 8.7555475e-07, -0.0021997013, 0.0003261454, 0.000113829214, 3.3664708e-06, -0.0023436933, 0.0002496961, 0.00011363622, 5.6730714e-06, -0.002449283, 0.00017273327, 0.00011166705, 7.769757e-06, -0.0025165125, 9.644509e-05, 0.00010803987, 9.6353915e-06, -0.0025460033, 2.1952763e-05, 0.00010289197, 1.1253385e-05, -0.002538917, -4.970307e-05, 9.637675e-05, 1.26117175e-05, -0.002496913, -0.00011757407, 8.8660614e-05, 1.3702878e-05, -0.0024220997, -0.00018081395, 7.9919846e-05, 1.4523757e-05, -0.0023169818, -0.00023868626, 7.0337504e-05, 1.50754695e-05, -0.002184403, -0.00029057014, 6.0100305e-05, 1.536312e-05, -0.0020274878, -0.00033596397, 4.9395687e-05, 1.5395543e-05, -0.0018495816, -0.00037448722, 3.8408944e-05, 1.518496e-05, -0.0016541894, -0.00040588036, 2.7320575e-05, 1.4746654e-05, -0.0014449162, -0.00043000278, 1.6303806e-05, 1.4098571e-05, -0.0012254084, -0.00044682936, 5.5223563e-06, 1.3260929e-05, -0.0009992969, -0.00045644512, -4.871546e-06, 1.2255797e-05, -0.0007701439, -0.00045903886, -1.4738881e-05, 1.1106677e-05, -0.00054139306, -0.0004548951, -2.3955274e-05, 9.838082e-06, -0.00031632345, -0.0004443856, -3.2412143e-05, 8.475117e-06, -9.800861e-05, -0.00042795928, -4.0017552e-05, 7.043077e-06, 0.00011071963, -0.00040613202, -4.669678e-05, 5.5670557e-06, 0.00030730182, -0.00037947576, -5.23926e-05, 4.0715845e-06, 0.00048947614, -0.00034860722, -5.706529e-05, 2.5802892e-06, 0.00065529795, -0.00031417652, -6.069237e-05, 1.1155827e-06, 0.0008031538, -0.0002768561, -6.326812e-05, -3.016111e-07, 0.00093176943, -0.00023732937, -6.480283e-05, -1.652098e-06, 0.001040213, -0.00019628023, -6.532189e-05, -2.9186162e-06, 0.0011278928, -0.00015438274, -6.486468e-05, -4.086e-06, 0.0011945489, -0.000112291564, -6.34833e-05, -5.141305e-06, 0.001240243, -7.0633265e-05, -6.124117e-05, -6.073893e-06, 0.0012653406, -2.9998188e-05, -5.821157e-05, -6.87548e-06, 0.0012704922, 9.066478e-06, -5.4476033e-05, -7.5401445e-06, 0.0012566097, 4.6062818e-05, -5.012275e-05, -8.064302e-06, 0.0012248404, 8.0547215e-05, -4.5244935e-05, -8.446648e-06, 0.0011765393, 0.00011213436, -3.9939183e-05, -8.688061e-06, 0.0011132385, 0.00014050014, -3.4303874e-05, -8.791489e-06, 0.0010366167, 0.00016538358, -2.8437618e-05, -8.761804e-06, 0.0009484669, 0.00018658763, -2.2437784e-05, -8.605636e-06, 0.00085066474, 0.00020397906, -1.639909e-05, -8.33119e-06, 0.00074513664, 0.00021748741, -1.0412333e-05, -7.948044e-06, 0.00063382904, 0.00022710294, -4.563222e-06, -7.4669465e-06, 0.0005186786, 0.00023287392, 1.0686539e-06, -6.8995923e-06, 0.000401584, 0.00023490313, 6.410718e-06, -6.2584086e-06, 0.00028437976, 0.0002333437, 1.1398149e-05, -5.55633e-06, 0.00016881226, 0.0002283944, 1.597447e-05, -4.8065845e-06, 5.6518104e-05, 0.00022029456, 2.0091995e-05, -4.0224795e-06, -5.0994746e-05, 0.00020931849, 2.3712108e-05, -3.2172018e-06, -0.00015236306, 0.0001957698, 2.680541e-05, -2.4036246e-06, -0.00024638147, 0.00017997542, 2.9351706e-05, -1.5941337e-06, -0.00033201274, 0.00016227973, 3.1339867e-05, -8.004638e-07, -0.00040839482, 0.00014303849, 3.2767566e-05, -3.3556752e-08, -0.00047484526, 0.00012261311, 3.3640874e-05, 6.9656414e-07, -0.0005308625, 0.00010136495, 3.397379e-05, 1.380899e-06, -0.0005761245, 7.965005e-05, 3.3787623e-05, 2.0115558e-06, -0.00061048503, 5.7814017e-05, 3.3110355e-05, 2.581815e-06, -0.0006339667, 3.6187455e-05, 3.197588e-05, 3.0861731e-06, -0.0006467532, 1.5081782e-05, 3.0423233e-05, 3.5203661e-06, -0.00064917805, -5.2144746e-06, 2.8495751e-05, 3.8813732e-06, -0.0006417128, -2.443884e-05, 2.624024e-05, 4.167402e-06, -0.00062495307, -4.2357522e-05, 2.3706087e-05, 4.3778564e-06, -0.0005996038, -5.8767506e-05, 2.0944432e-05, 4.5132883e-06, -0.0005664634, -7.349806e-05, 1.8007306e-05, 4.5753336e-06, -0.00052640727, -8.641171e-05, 1.4946819e-05, 4.5666357e-06, -0.00048037132, -9.7404685e-05, 1.1814389e-05, 4.490758e-06, -0.00042933473, -0.00010640679, 8.6600085e-06, 4.3520886e-06, -0.00037430358, -0.000113380855, 5.5315704e-06, 4.155732e-06, -0.0003162945, -0.00011832167, 2.4742617e-06, 3.907401e-06, -0.00025631895, -0.000121254496, -4.6997877e-07, 3.613304e-06, -0.00019536859, -0.00012223326, -3.2629237e-06, 3.2800256e-06, -0.00013440137, -0.00012133831, -5.870446e-06, 2.914413e-06, -7.432899e-05, -0.000118673976, -8.262828e-06, 2.5234622e-06, -1.600553e-05, -0.00011436584, -1.0414987e-05, 2.1142048e-06, 3.9782444e-05, -0.00010855784, -1.2306627e-05, 1.6936041e-06, 9.232428e-05, -0.00010140926, -1.3922302e-05, 1.2684541e-06, 0.00014099214, -9.309159e-05, -1.5251419e-05, 8.45287e-07, 0.00018524638, -8.378541e-05, -1.6288155e-05, 4.302888e-07, 0.00022463918, -7.3677234e-05, -1.7031312e-05, 2.9224458e-08, 0.0002588169, -6.29565e-05, -1.7484113e-05, -3.5262744e-07, 0.0002875207, -5.1812534e-05, -1.7653942e-05, -7.105295e-07, 0.0003105858, -4.043184e-05, -1.7552025e-05, -1.0403297e-06, 0.00032793934, -2.8995384e-05, -1.7193088e-05, -1.3384947e-06, 0.0003395971, -1.7676197e-05, -1.659496e-05, -1.6021322e-06, 0.000345659, -6.6371917e-06, -1.5778161e-05, -1.8290033e-06, 0.0003463033, 3.970771e-06, -1.4765471e-05, -2.0175235e-06, 0.0003417805, 1.40105485e-05, -1.3581472e-05, -2.166755e-06, 0.00033240582, 2.3360086e-05, -1.2252103e-05, -2.2763893e-06, 0.00031855155, 3.1913507e-05, -1.08042095e-05, -2.3467212e-06, 0.0003006387, 3.9581897e-05, -9.265097e-06, -2.378615e-06, 0.00027912838, 4.6293808e-05, -7.662104e-06, -2.3734647e-06, 0.00025451303, 5.1995485e-05, -6.022192e-06, -2.333147e-06, 0.00022730745, 5.6650795e-05, -4.3715686e-06, -2.2599704e-06, 0.0001980403, 6.0240916e-05, -2.7353294e-06, -2.15662e-06, 0.00016724532, 6.276379e-05, -1.1371408e-06, -2.0260989e-06, 0.0001354533, 6.4233325e-05, 4.010435e-07, -1.8716687e-06, 0.00010318427, 6.467843e-05, 1.8592249e-06, -1.6967887e-06, 7.094028e-05, 6.414185e-05, 3.2195635e-06, -1.5050541e-06, 3.9198825e-05, 6.267888e-05, 4.466538e-06, -1.3001369e-06, 8.406919e-06, 6.035591e-05, 5.587065e-06, -1.0857268e-06, -2.1024085e-05, 5.7248908e-05, 6.570575e-06, -8.65476e-07, -4.872289e-05, 5.3441847e-05, 7.409048e-06, -6.4294665e-07, -7.436183e-05, 4.9025046e-05, 8.097009e-06, -4.2156222e-07, -9.765966e-05, 4.4093536e-05, 8.631489e-06, -2.0456325e-07, -0.00011838346, 3.874541e-05, 9.011942e-06, 5.031821e-09, -0.0001363498, 3.3080214e-05, 9.240142e-06, 2.0446087e-07, -0.00015142508, 2.7197406e-05, 9.320041e-06, 3.9124672e-07, -0.00016352505, 2.1194879e-05, 9.257604e-06, 5.6322017e-07, -0.00017261377, 1.51675795e-05, 9.060629e-06, 7.185373e-07, -0.00017870174, 9.2062355e-06, 8.738533e-06, 8.5569127e-07, -0.00018184353, 3.3962156e-06, 8.302143e-06, 9.735182e-07, -0.00018213484, -2.1834817e-06, 7.7634595e-06, 1.0711982e-06, -0.00017970912, -7.4610953e-06, 7.135425e-06, 1.1482504e-06, -0.00017473368, -1.237282e-05, 6.4316873e-06, 1.2045243e-06, -0.00016740568, -1.6863367e-05, 5.666358e-06, 1.2401855e-06, -0.00015794765, -2.0886377e-05, 4.853784e-06, 1.2556984e-06, -0.00014660307, -2.440468e-05, 4.0083223e-06, 1.2518045e-06, -0.00013363162, -2.7390399e-05, 3.1441236e-06, 1.229498e-06, -0.00011930462, -2.9824914e-05, 2.2749355e-06, 1.1899991e-06, -0.00010390044, -3.1698703e-05, 1.4139143e-06, 1.1347245e-06, -8.769998e-05, -3.301103e-05, 5.734608e-07, 1.065257e-06, -7.0982365e-05, -3.376954e-05, -2.3493e-07, 9.833144e-07, -5.4020962e-05, -3.398973e-05, -1.0007943e-06, 8.9071654e-07, -3.7079502e-05, -3.3694363e-05, -1.714806e-06, 7.893539e-07, -2.0408694e-05, -3.2912747e-05, -2.3688601e-06, 6.811561e-07, -4.24309e-06, -3.168001e-05, -2.9561345e-06, 5.6806107e-07, 1.1201599e-05, -3.003628e-05, -3.4711288e-06, 4.519859e-07, 2.5730804e-05, -2.8025852e-05, -3.9096826e-06, 3.3479944e-07, 3.917297e-05, -2.569633e-05, -4.268973e-06, 2.1829676e-07, 5.1380986e-05, -2.3097758e-05, -4.547491e-06, 1.041761e-07, 6.223319e-05, -2.0281763e-05, -4.7450003e-06, -5.981753e-09, 7.163397e-05, -1.7300701e-05, -4.862482e-06, -1.107313e-07, 7.9513884e-05, -1.4206852e-05, -4.902057e-06, -2.0877722e-07, 8.5829444e-05, -1.1051647e-05, -4.8669017e-06, -2.9898644e-07, 9.0562535e-05, -7.884938e-06, -4.761151e-06, -3.8039704e-07, 9.371941e-05, -4.754341e-06, -4.589788e-06, -4.5222438e-07, 9.532947e-05, -1.7046308e-06, -4.35853e-06, -5.1386417e-07, 9.5443655e-05, 1.2227831e-06, -4.073709e-06, -5.648927e-07, 9.413267e-05, 3.990312e-06, -3.7421453e-06, -6.050644e-07, 9.148501e-05, 6.5645604e-06, -3.3710255e-06, -6.3430696e-07, 8.760472e-05, 8.916621e-06, -2.9677767e-06, -6.52714e-07, 8.260916e-05, 1.1022283e-05, -2.539944e-06, -6.605356e-07, 7.662656e-05, 1.2862173e-05, -2.0950731e-06, -6.581671e-07, 6.9793634e-05, 1.4421801e-05, -1.6405986e-06, -6.461362e-07, 6.2253115e-05, 1.5691545e-05, -1.183738e-06, -6.250886e-07, 5.4151365e-05, 1.6666554e-05, -7.313957e-07, -5.957729e-07, 4.563598e-05, 1.7346594e-05, -2.900748e-07, -5.590244e-07, 3.6853584e-05, 1.7735827e-05, 1.3419942e-07, -5.157483e-07, 2.794767e-05, 1.7842533e-05, 5.359465e-07, -4.6690323e-07, 1.9056624e-05, 1.767879e-05, 9.102856e-07, -4.1348426e-07, 1.0311924e-05, 1.726012e-05, 1.2529792e-06, -3.5650626e-07, 1.836507e-06, 1.660507e-05, 1.5604652e-06, -2.9698796e-07, -6.2566364e-06, 1.5734817e-05, 1.8298765e-06, -2.3593658e-07, -1.3865663e-05, 1.4672701e-05, 2.0590508e-06, -1.7433346e-07, -2.0900854e-05, 1.3443791e-05, 2.246528e-06, -1.13120706e-07, -2.7285358e-05, 1.20744235e-05, 2.391539e-06, -5.318905e-08, -3.295571e-05, 1.0591746e-05, 2.4939823e-06, 4.6328443e-09, -3.786214e-05, 9.02328e-06, 2.5543943e-06, 5.9587748e-08, -4.1968633e-05, 7.396488e-06, 2.5739098e-06, 1.1099764e-07, -4.5252804e-05, 5.738375e-06, 2.554217e-06, 1.5826997e-07, -4.7705584e-05, 4.0751033e-06, 2.497505e-06, 2.009023e-07, -4.9330694e-05, 2.4316482e-06, 2.406407e-06, 2.3848548e-07, -5.0143983e-05, 8.314821e-07, 2.2839404e-06, 2.7070516e-07, -5.01726e-05, -7.037013e-07, 2.1334424e-06, 2.973419e-07, -4.9454047e-05, -2.1542228e-06, 1.9585061e-06, 3.1826983e-07, -4.8035115e-05, -3.502613e-06, 1.7629134e-06, 3.3345404e-07, -4.597075e-05, -4.733766e-06, 1.5505706e-06, 3.4294666e-07, -4.3322838e-05, -5.835049e-06, 1.3254444e-06, 3.4688188e-07, -4.015894e-05, -6.7963683e-06, 1.091499e-06, 3.4546997e-07, -3.655102e-05, -7.6102024e-06, 8.526388e-07, 3.3899056e-07, -3.2574175e-05, -8.271582e-06, 6.126518e-07, 3.2778505e-07, -2.8305343e-05, -8.778047e-06, 3.751598e-07, 3.1224855e-07, -2.3822091e-05, -9.129557e-06, 1.435725e-07, 2.9282148e-07, -1.9201418e-05, -9.328378e-06, -7.8953136e-08, 2.6998077e-07, -1.4518649e-05, -9.378936e-06, -2.895475e-07, 2.44231e-07, -9.846386e-06, -9.287646e-06, -4.856571e-07, 2.160956e-07, -5.2535684e-06, -9.062723e-06, -6.650671e-07, 1.8610817e-07, -8.0462104e-07, -8.713968e-06, -8.259181e-07, 1.5480401e-07, 3.4412838e-06, -8.252551e-06, -9.667165e-07, 1.2271214e-07, 7.4308523e-06, -7.690779e-06, -1.0863387e-06, 9.034764e-08, 1.1117177e-05, -7.04185e-06, -1.1840305e-06, 5.820481e-08, 1.4460125e-05, -6.3196244e-06, -1.2593999e-06, 2.6750717e-08, 1.7426608e-05, -5.5383794e-06, -1.312406e-06, -3.5803926e-09, 1.999073e-05, -4.71258e-06, -1.3433419e-06, -3.2391956e-08, 2.213383e-05, -3.8566545e-06, -1.3528147e-06, -5.932917e-08, 2.3844408e-05, -2.984781e-06, -1.3417213e-06, -8.408225e-08, 2.5117946e-05, -2.1106891e-06, -1.3112208e-06, -1.0638886e-07, 2.595664e-05, -1.2474783e-06, -1.2627047e-06, -1.2603569e-07, 2.6369045e-05, -4.0745232e-07, -1.1977652e-06, -1.4285932e-07, 2.6369638e-05, 3.980239e-07, -1.1181614e-06, -1.5674614e-07, 2.5978317e-05, 1.1586486e-06, -1.0257855e-06, -1.6763174e-07, 2.521984e-05, 1.8652848e-06, -9.2262803e-07, -1.754994e-07, 2.4123232e-05, 2.5100396e-06, -8.1074336e-07, -1.8037807e-07, 2.2721133e-05, 3.0863212e-06, -6.9221653e-07, -1.8233975e-07, 2.104915e-05, 3.5888745e-06, -5.691303e-07, -1.8149628e-07, 1.9145182e-05, 4.0137943e-06, -4.4353462e-07, -1.7799583e-07, 1.7048738e-05, 4.358518e-06, -3.174176e-07, -1.7201887e-07, 1.4800284e-05, 4.6217983e-06, -1.92679e-07, -1.6377396e-07, 1.2440583e-05, 4.80366e-06, -7.1106214e-08, -1.5349329e-07, 1.0010085e-05, 4.9053356e-06, 4.564679e-08, -1.414281e-07, 7.5483367e-06, 4.9291907e-06, 1.5607766e-07, -1.2784398e-07, 5.0934354e-06, 4.8786324e-06, 2.5885066e-07, -1.1301628e-07, 2.6815364e-06, 4.75801e-06, 3.5280843e-07, -9.7225495e-08, 3.4640763e-07, 4.5725033e-06, 4.3698057e-07, -8.075291e-08, -1.8809568e-06, 4.328006e-06, 5.1058913e-07, -6.3876314e-08, -3.9726624e-06, 4.031004e-06, 5.730506e-07, -4.68661e-08, -5.9041804e-06, 3.6884505e-06, 6.239756e-07, -2.9981543e-08, -7.654547e-06, 3.3076383e-06, 6.631648e-07, -1.3467543e-08, -9.206506e-06, 2.8960771e-06, 6.906032e-07, 2.448364e-09, -1.0546583e-05, 2.4613707e-06, 7.06451e-07, 1.7558524e-08, -1.1665106e-05, 2.011099e-06, 7.1103284e-07, 3.16773e-08, -1.2556163e-05, 1.5527066e-06, 7.048254e-07, 4.4642764e-08, -1.32175055e-05, 1.0933995e-06, 6.884425e-07, 5.6317965e-08, -1.3650413e-05, 6.400486e-07, 6.626196e-07, 6.659174e-08, -1.3859495e-05, 1.9910387e-07, 6.2819674e-07, 7.5379134e-08, -1.3852466e-05, -2.2348063e-07, 5.861014e-07, 8.26214e-08, -1.36398785e-05, -6.223117e-07, 5.3733015e-07, 8.828558e-08, -1.3234832e-05, -9.926099e-07, 4.8293055e-07, 9.236379e-08, -1.2652653e-05, -1.3302508e-06, 4.2398335e-07, 9.487207e-08, -1.1910556e-05, -1.6317953e-06, 3.6158445e-07, 9.584904e-08, -1.1027305e-05, -1.8945062e-06, 2.968282e-07, 9.535421e-08, -1.0022853e-05, -2.1163567e-06, 2.3079103e-07, 9.3466085e-08, -8.917988e-06, -2.2960246e-06, 1.6451636e-07, 9.028008e-08, -7.733988e-06, -2.432879e-06, 9.9000744e-08, 8.59063e-08, -6.4922774e-06, -2.5269558e-06, 3.5181213e-08, 8.046717e-08, -5.214102e-06, -2.5789248e-06, -2.607566e-08, 7.4095034e-08, -3.920223e-06, -2.5900495e-06, -8.398331e-08, 6.6929715e-08, -2.6306316e-06, -2.5621393e-06, -1.3784297e-07, 5.9116044e-08, -1.3642878e-06, -2.497496e-06, -1.8704985e-07, 5.080151e-08, -1.3889007e-07, -2.3988569e-06, -2.3109749e-07, 4.2133905e-08, 1.0293274e-06, -2.2693312e-06, -2.6958065e-07, 3.325912e-08, 2.1257656e-06, -2.1123374e-06, -3.021964e-07, 2.4319084e-08, 3.1375978e-06, -1.9315373e-06, -3.2874362e-07, 1.5449821e-08, 4.0538753e-06, -1.7307689e-06, -3.491211e-07, 6.779738e-09, 4.8655984e-06, -1.5139818e-06, -3.6332432e-07, -1.5719323e-09, 5.565757e-06, -1.2851727e-06, -3.7144062e-07, -9.496452e-09, 6.149339e-06, -1.0483236e-06, -3.7364367e-07, -1.689669e-08, 6.6133052e-06, -8.0734367e-07, -3.7018663e-07, -2.3688003e-08, 6.956543e-06, -5.660143e-07, -3.6139448e-07, -2.9798889e-08, 7.1797876e-06, -3.2793946e-07, -3.476559e-07, -3.5171418e-08, 7.285522e-06, -9.650032e-08, -3.294142e-07, -3.976144e-08, 7.2778557e-06, 1.2518392e-07, -3.0715825e-07, -4.3538552e-08, 7.162385e-06, 3.342899e-07, -2.814129e-07, -4.648593e-08, 6.9460384e-06, 5.283177e-07, -2.527295e-07, -4.859987e-08, 6.636909e-06, 7.051124e-07, -2.2167647e-07, -4.9889252e-08, 6.244076e-06, 8.628794e-07, -1.8882989e-07, -5.0374776e-08, 5.7774255e-06, 1.0001936e-06, -1.5476468e-07, -5.0088094e-08, 5.247463e-06, 1.116003e-06, -1.200461e-07, -4.907079e-08, 4.6651253e-06, 1.2096259e-06, -8.522175e-08, -4.7373316e-08, 4.041601e-06, 1.2807433e-06, -5.081436e-08, -4.5053785e-08, 3.3881486e-06, 1.3293862e-06, -1.7315188e-08, -4.2176744e-08, 2.7159272e-06, 1.3559182e-06, 1.4821778e-08, -3.8811912e-08, 2.0358364e-06, 1.361014e-06, 4.5184727e-08, -3.5032883e-08, 1.3583644e-06, 1.3456342e-06, 7.340813e-08, -3.0915857e-08, 6.9345475e-07, 1.3109972e-06, 9.917594e-08, -2.6538357e-08, 5.038252e-08, 1.2585489e-06, 1.2222388e-07, -2.197805e-08, -5.6234967e-07, 1.1899299e-06, 1.4234087e-07, -1.731155e-08, -1.1371013e-06, 1.106942e-06, 1.5936959e-07, -1.2613351e-08, -1.6671659e-06, 1.0115133e-06, 1.7320627e-07, -7.954819e-09, -2.1468254e-06, 9.0566357e-07, 1.8379957e-07, -3.4032754e-09, -2.571387e-06, 7.9147003e-07, 1.9114884e-07, 9.788003e-10, -2.9372043e-06, 6.710333e-07, 1.9530167e-07, 5.134469e-09, -3.2416801e-06, 5.464454e-07, 1.9635088e-07, 9.0129095e-09, -3.4832542e-06, 4.1975866e-07, 1.9443092e-07, 1.2569879e-08, -3.6613771e-06, 2.9295762e-07, 1.8971389e-07, 1.576805e-08, -3.776469e-06, 1.6793253e-07, 1.8240512e-07, 1.8577236e-08, -3.8298663e-06, 4.6455742e-08, 1.7273852e-07, 2.0974484e-08, -3.823758e-06, -6.983869e-08, 1.609718e-07, 2.2944084e-08, -3.7611119e-06, -1.794728e-07, 1.4738134e-07, 2.4477433e-08, -3.6455922e-06, -2.8113908e-07, 1.3225736e-07, 2.5572833e-08, -3.4814725e-06, -3.737116e-07, 1.1589875e-07, 2.6235176e-08, -3.273541e-06, -4.562541e-07, 9.860837e-08, 2.6475552e-08, -3.0270073e-06, -5.280246e-07, 8.068825e-08, 2.6310792e-08, -2.7474011e-06, -5.884772e-07, 6.243519e-08, 2.5762928e-08, -2.4404778e-06, -6.372605e-07, 4.4136584e-08, 2.4858627e-08, -2.1121195e-06, -6.7421354e-07, 2.6066619e-08, 2.3628562e-08, -1.768243e-06, -6.993591e-07, 8.482815e-09, 2.2106766e-08, -1.4147099e-06, -7.1289423e-07, -8.376974e-09, 2.032996e-08, -1.0572415e-06, -7.1517906e-07, -2.429716e-08, 1.8336882e-08, -7.013413e-07, -7.0672354e-07, -3.908654e-08, 1.6167615e-08, -3.522233e-07, -6.881726e-07, -5.2579967e-08, 1.3862916e-08, -1.4748624e-08, -6.6029e-07, -6.4639536e-08, 1.146359e-08, 3.066297e-07, -6.239414e-07, -7.515533e-08, 9.009873e-09, 6.079131e-07, -5.800763e-07, -8.4045666e-08, 6.5408656e-09, 8.85595e-07, -5.2971006e-07, -9.125701e-08, 4.0940042e-09, 1.1366892e-06, -4.7390563e-07, -9.676333e-08, 1.7045872e-09, 1.3587492e-06, -4.1375532e-07, -1.0056523e-07, -5.946482e-10, 1.5498778e-06, -3.5036328e-07, -1.02688595e-07, -2.7738878e-09, 1.7087299e-06, -2.8482845e-07, -1.0318301e-07, -4.806542e-09, 1.8345047e-06, -2.1822848e-07, -1.021199e-07, -6.669485e-09, 1.926932e-06, -1.5160478e-07, -9.959034e-08, -8.343233e-09, 1.9862505e-06, -8.594872e-08, -9.570284e-08, -9.812055e-09, 2.0131788e-06, -2.2189392e-08, -9.058082e-08, -1.1064026e-08, 2.0088828e-06, 3.881723e-08, -8.43601e-08, -1.2091022e-08, 1.9749357e-06, 9.629747e-08, -7.718627e-08, -1.2888656e-08, 1.913276e-06, 1.4956747e-07, -6.921202e-08, -1.345616e-08, 1.8261597e-06, 1.98039e-07, -6.059457e-08, -1.3796225e-08, 1.7161124e-06, 2.4122363e-07, -5.149311e-08, -1.3914792e-08, 1.5858784e-06, 2.7873506e-07, -4.206631e-08, -1.3820808e-08, 1.4383693e-06, 3.1029006e-07, -3.2470016e-08, -1.3525944e-08, 1.2766128e-06, 3.3570754e-07, -2.2855051e-08, -1.3044296e-08, 1.103702e-06, 3.549065e-07, -1.336523e-08, -1.2392054e-08, 9.2274604e-07, 3.6790215e-07, -4.135552e-09, -1.1587158e-08, 7.3682355e-07, 3.748013e-07, 4.709376e-09, -1.0648952e-08, 5.489381e-07, 3.757961e-07, 1.3056691e-08, -9.5978265e-09, 3.619772e-07, 3.7115723e-07, 2.080638e-08, -8.454863e-09, 1.7867491e-07, 3.6122603e-07, 2.7872154e-08, -7.24149e-09, 1.5789132e-09, 3.4640595e-07, 3.418205e-08, -5.979147e-09, -1.6697864e-07, 3.2715363e-07, 3.9678834e-08, -4.688963e-09, -3.2490524e-07, 3.039695e-07, 4.4320114e-08, -3.391461e-09, -4.7036752e-07, 2.7738824e-07, 4.8078263e-08, -2.1062794e-09, -6.0180605e-07, 2.4796915e-07, 5.0940116e-08, -8.5192514e-10, -7.1794517e-07, 2.1628675e-07, 5.2906476e-08, 3.5444864e-10, -8.1779837e-07, 1.8292133e-07, 5.3991403e-08, 1.4972308e-09, -9.0066885e-07, 1.4845017e-07, 5.4221392e-08, 2.5625104e-09, -9.66146e-07, 1.134391e-07, 5.363435e-08, 3.5382006e-09, -1.0140974e-06, 7.8434596e-08, 5.227851e-08, 4.414131e-09, -1.0446577e-06, 4.3956618e-08, 5.0211185e-08, 5.182105e-09, -1.0582135e-06, 1.0492179e-08, 4.7497505e-08, 5.8359273e-09, -1.0553852e-06, -2.1510338e-08, 4.420905e-08, 6.371399e-09, -1.0370072e-06, -5.1645944e-08, 4.0422485e-08, 6.7862826e-09, -1.0041043e-06, -7.955698e-08, 3.621818e-08, 7.080242e-09, -9.578679e-07, -1.04936156e-07, 3.167881e-08, 7.254754e-09, -8.9962964e-07, -1.2752865e-07, 2.688805e-08, 7.3129995e-09};
endpackage
`endif
