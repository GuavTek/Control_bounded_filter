`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam N = 4;
	localparam M = 4;
	localparam real Lfr[0:3] = {0.9933908, 0.9933908, 0.9848978, 0.9848978};
	localparam real Lfi[0:3] = {0.030115983, -0.030115983, 0.012144258, -0.012144258};
	localparam real Lbr[0:3] = {0.9933908, 0.9933908, 0.9848978, 0.9848978};
	localparam real Lbi[0:3] = {0.030115983, -0.030115983, 0.012144258, -0.012144258};
	localparam real Wfr[0:3] = {2.0204313e-06, 2.0204313e-06, 6.0135073e-07, 6.0135073e-07};
	localparam real Wfi[0:3] = {7.631857e-08, -7.631857e-08, 1.1569381e-06, -1.1569381e-06};
	localparam real Wbr[0:3] = {-2.0204313e-06, -2.0204313e-06, -6.0135073e-07, -6.0135073e-07};
	localparam real Wbi[0:3] = {-7.631857e-08, 7.631857e-08, -1.1569381e-06, 1.1569381e-06};
	localparam real Ffr[0:3][0:99] = '{
		'{743.8243, 45.974236, -3.1845877, 0.020513162, 766.31213, 43.9743, -3.1971812, 0.024781875, 787.7957, 41.9571, -3.206581, 0.028974663, 808.2667, 39.924755, -3.2128172, 0.033088468, 827.71826, 37.87939, -3.2159226, 0.037120353, 846.1443, 35.82311, -3.2159326, 0.041067485, 863.5399, 33.757996, -3.2128851, 0.044927154, 879.9012, 31.686125, -3.206821, 0.048696768, 895.2252, 29.609549, -3.1977825, 0.052373838, 909.51025, 27.530298, -3.1858149, 0.05595601, 922.75543, 25.450384, -3.1709654, 0.059441045, 934.9609, 23.371792, -3.1532838, 0.06282682, 946.12775, 21.296482, -3.1328213, 0.066111326, 956.25824, 19.226383, -3.1096315, 0.069292694, 965.35535, 17.163404, -3.0837703, 0.07236916, 973.42316, 15.109415, -3.0552945, 0.07533909, 980.46655, 13.066261, -3.0242636, 0.07820096, 986.4915, 11.03575, -2.9907384, 0.08095338, 991.5047, 9.019657, -2.9547813, 0.083595075, 995.51385, 7.0197234, -2.9164562, 0.0861249, 998.5274, 5.0376506, -2.8758287, 0.088541806, 1000.55475, 3.075104, -2.8329659, 0.090844885, 1001.606, 1.1337103, -2.7879357, 0.09303336, 1001.69226, -0.7849449, -2.7408075, 0.09510654, 1000.82513, -2.6793163, -2.691652, 0.09706387},
		'{743.8243, 45.974236, -3.1845877, 0.020513162, 766.31213, 43.9743, -3.1971812, 0.024781875, 787.7957, 41.9571, -3.206581, 0.028974663, 808.2667, 39.924755, -3.2128172, 0.033088468, 827.71826, 37.87939, -3.2159226, 0.037120353, 846.1443, 35.82311, -3.2159326, 0.041067485, 863.5399, 33.757996, -3.2128851, 0.044927154, 879.9012, 31.686125, -3.206821, 0.048696768, 895.2252, 29.609549, -3.1977825, 0.052373838, 909.51025, 27.530298, -3.1858149, 0.05595601, 922.75543, 25.450384, -3.1709654, 0.059441045, 934.9609, 23.371792, -3.1532838, 0.06282682, 946.12775, 21.296482, -3.1328213, 0.066111326, 956.25824, 19.226383, -3.1096315, 0.069292694, 965.35535, 17.163404, -3.0837703, 0.07236916, 973.42316, 15.109415, -3.0552945, 0.07533909, 980.46655, 13.066261, -3.0242636, 0.07820096, 986.4915, 11.03575, -2.9907384, 0.08095338, 991.5047, 9.019657, -2.9547813, 0.083595075, 995.51385, 7.0197234, -2.9164562, 0.0861249, 998.5274, 5.0376506, -2.8758287, 0.088541806, 1000.55475, 3.075104, -2.8329659, 0.090844885, 1001.606, 1.1337103, -2.7879357, 0.09303336, 1001.69226, -0.7849449, -2.7408075, 0.09510654, 1000.82513, -2.6793163, -2.691652, 0.09706387},
		'{741.83435, 45.861446, -3.1145601, 0.2656197, 764.2799, 43.927692, -3.0076368, 0.25940147, 785.7689, 42.035126, -2.9027734, 0.2532713, 806.32184, 40.183224, -2.7999477, 0.24722889, 825.95886, 38.371468, -2.699138, 0.24127385, 844.6999, 36.59935, -2.6003213, 0.23540583, 862.5647, 34.86634, -2.5034757, 0.22962445, 879.5727, 33.171936, -2.4085786, 0.22392929, 895.743, 31.515614, -2.3156075, 0.2183199, 911.09454, 29.89686, -2.2245402, 0.21279582, 925.646, 28.315166, -2.1353538, 0.20735663, 939.41583, 26.770018, -2.0480258, 0.2020018, 952.42206, 25.260904, -1.9625337, 0.19673084, 964.6826, 23.787321, -1.8788545, 0.1915432, 976.2152, 22.348759, -1.7969657, 0.18643838, 987.0372, 20.944714, -1.7168448, 0.18141583, 997.1656, 19.574684, -1.638469, 0.17647494, 1006.61743, 18.238169, -1.5618157, 0.17161517, 1015.40924, 16.934671, -1.4868623, 0.16683589, 1023.5575, 15.663694, -1.4135864, 0.16213652, 1031.0782, 14.424747, -1.3419652, 0.15751645, 1037.9875, 13.21734, -1.2719765, 0.15297502, 1044.3008, 12.040984, -1.2035977, 0.14851162, 1050.0336, 10.895195, -1.1368065, 0.14412557, 1055.201, 9.779492, -1.0715808, 0.13981622},
		'{741.83435, 45.861446, -3.1145601, 0.2656197, 764.2799, 43.927692, -3.0076368, 0.25940147, 785.7689, 42.035126, -2.9027734, 0.2532713, 806.32184, 40.183224, -2.7999477, 0.24722889, 825.95886, 38.371468, -2.699138, 0.24127385, 844.6999, 36.59935, -2.6003213, 0.23540583, 862.5647, 34.86634, -2.5034757, 0.22962445, 879.5727, 33.171936, -2.4085786, 0.22392929, 895.743, 31.515614, -2.3156075, 0.2183199, 911.09454, 29.89686, -2.2245402, 0.21279582, 925.646, 28.315166, -2.1353538, 0.20735663, 939.41583, 26.770018, -2.0480258, 0.2020018, 952.42206, 25.260904, -1.9625337, 0.19673084, 964.6826, 23.787321, -1.8788545, 0.1915432, 976.2152, 22.348759, -1.7969657, 0.18643838, 987.0372, 20.944714, -1.7168448, 0.18141583, 997.1656, 19.574684, -1.638469, 0.17647494, 1006.61743, 18.238169, -1.5618157, 0.17161517, 1015.40924, 16.934671, -1.4868623, 0.16683589, 1023.5575, 15.663694, -1.4135864, 0.16213652, 1031.0782, 14.424747, -1.3419652, 0.15751645, 1037.9875, 13.21734, -1.2719765, 0.15297502, 1044.3008, 12.040984, -1.2035977, 0.14851162, 1050.0336, 10.895195, -1.1368065, 0.14412557, 1055.201, 9.779492, -1.0715808, 0.13981622}};
	localparam real Ffi[0:3][0:99] = '{
		'{-909.9477, 56.318283, 1.1170552, -0.14624423, -881.5327, 57.330624, 1.0137653, -0.1446599, -852.62823, 58.276043, 0.91077894, -0.1429575, -823.2678, 59.154465, 0.8081901, -0.14114006, -793.4849, 59.965878, 0.70609146, -0.13921075, -763.3131, 60.710327, 0.6045741, -0.13717276, -732.78577, 61.387928, 0.5037274, -0.13502938, -701.9363, 61.99886, 0.40363896, -0.1327839, -670.798, 62.543354, 0.3043947, -0.13043976, -639.40393, 63.021717, 0.20607851, -0.12800038, -607.78723, 63.434296, 0.10877256, -0.12546922, -575.9805, 63.78151, 0.0125569245, -0.12284985, -544.01654, 64.06383, -0.0824903, -0.12014582, -511.92746, 64.281784, -0.1762931, -0.11736075, -479.74536, 64.43596, -0.26877755, -0.11449827, -447.502, 64.52698, -0.35987192, -0.111562066, -415.22882, 64.55554, -0.44950667, -0.108555816, -382.95676, 64.522385, -0.53761446, -0.10548326, -350.71658, 64.4283, -0.6241303, -0.102348104, -318.53848, 64.27412, -0.70899147, -0.09915412, -286.45233, 64.06072, -0.79213756, -0.09590506, -254.48747, 63.789047, -0.87351054, -0.09260468, -222.67284, 63.460064, -0.9530549, -0.089256756, -191.03679, 63.074787, -1.0307175, -0.08586505, -159.60725, 62.634277, -1.1064473, -0.08243332},
		'{909.9477, -56.318283, -1.1170552, 0.14624423, 881.5327, -57.330624, -1.0137653, 0.1446599, 852.62823, -58.276043, -0.91077894, 0.1429575, 823.2678, -59.154465, -0.8081901, 0.14114006, 793.4849, -59.965878, -0.70609146, 0.13921075, 763.3131, -60.710327, -0.6045741, 0.13717276, 732.78577, -61.387928, -0.5037274, 0.13502938, 701.9363, -61.99886, -0.40363896, 0.1327839, 670.798, -62.543354, -0.3043947, 0.13043976, 639.40393, -63.021717, -0.20607851, 0.12800038, 607.78723, -63.434296, -0.10877256, 0.12546922, 575.9805, -63.78151, -0.0125569245, 0.12284985, 544.01654, -64.06383, 0.0824903, 0.12014582, 511.92746, -64.281784, 0.1762931, 0.11736075, 479.74536, -64.43596, 0.26877755, 0.11449827, 447.502, -64.52698, 0.35987192, 0.111562066, 415.22882, -64.55554, 0.44950667, 0.108555816, 382.95676, -64.522385, 0.53761446, 0.10548326, 350.71658, -64.4283, 0.6241303, 0.102348104, 318.53848, -64.27412, 0.70899147, 0.09915412, 286.45233, -64.06072, 0.79213756, 0.09590506, 254.48747, -63.789047, 0.87351054, 0.09260468, 222.67284, -63.460064, 0.9530549, 0.089256756, 191.03679, -63.074787, 1.0307175, 0.08586505, 159.60725, -62.634277, 1.1064473, 0.08243332},
		'{-2770.766, 102.199974, -4.9312606, 0.18171343, -2719.9124, 101.213486, -4.894612, 0.1821949, -2669.554, 100.21841, -4.857218, 0.1825936, -2619.6953, 99.21537, -4.819115, 0.18291183, -2570.3398, 98.204994, -4.780339, 0.18315186, -2521.4915, 97.187874, -4.7409244, 0.18331595, -2473.153, 96.1646, -4.700905, 0.18340631, -2425.328, 95.13572, -4.6603136, 0.18342508, -2378.018, 94.10181, -4.619183, 0.1833744, -2331.2268, 93.0634, -4.577544, 0.18325639, -2284.9553, 92.02101, -4.5354285, 0.18307306, -2239.2063, 90.97515, -4.492866, 0.18282644, -2193.9807, 89.92633, -4.4498854, 0.18251851, -2149.2803, 88.875015, -4.4065156, 0.18215123, -2105.1062, 87.821686, -4.362785, 0.1817265, -2061.459, 86.76679, -4.31872, 0.18124618, -2018.3395, 85.710785, -4.274348, 0.18071212, -1975.7483, 84.654076, -4.2296934, 0.18012613, -1933.6854, 83.59711, -4.184783, 0.17948996, -1892.1511, 82.54026, -4.1396403, 0.17880537, -1851.1451, 81.48395, -4.0942893, 0.17807403, -1810.667, 80.428535, -4.0487537, 0.17729764, -1770.7163, 79.3744, -4.0030556, 0.17647782, -1731.2924, 78.3219, -3.9572175, 0.17561617, -1692.3942, 77.27138, -3.9112604, 0.17471428},
		'{2770.766, -102.199974, 4.9312606, -0.18171343, 2719.9124, -101.213486, 4.894612, -0.1821949, 2669.554, -100.21841, 4.857218, -0.1825936, 2619.6953, -99.21537, 4.819115, -0.18291183, 2570.3398, -98.204994, 4.780339, -0.18315186, 2521.4915, -97.187874, 4.7409244, -0.18331595, 2473.153, -96.1646, 4.700905, -0.18340631, 2425.328, -95.13572, 4.6603136, -0.18342508, 2378.018, -94.10181, 4.619183, -0.1833744, 2331.2268, -93.0634, 4.577544, -0.18325639, 2284.9553, -92.02101, 4.5354285, -0.18307306, 2239.2063, -90.97515, 4.492866, -0.18282644, 2193.9807, -89.92633, 4.4498854, -0.18251851, 2149.2803, -88.875015, 4.4065156, -0.18215123, 2105.1062, -87.821686, 4.362785, -0.1817265, 2061.459, -86.76679, 4.31872, -0.18124618, 2018.3395, -85.710785, 4.274348, -0.18071212, 1975.7483, -84.654076, 4.2296934, -0.18012613, 1933.6854, -83.59711, 4.184783, -0.17948996, 1892.1511, -82.54026, 4.1396403, -0.17880537, 1851.1451, -81.48395, 4.0942893, -0.17807403, 1810.667, -80.428535, 4.0487537, -0.17729764, 1770.7163, -79.3744, 4.0030556, -0.17647782, 1731.2924, -78.3219, 3.9572175, -0.17561617, 1692.3942, -77.27138, 3.9112604, -0.17471428}};
	localparam real Fbr[0:3][0:99] = '{
		'{-743.8243, 45.974236, 3.1845877, 0.020513162, -766.31213, 43.9743, 3.1971812, 0.024781875, -787.7957, 41.9571, 3.206581, 0.028974663, -808.2667, 39.924755, 3.2128172, 0.033088468, -827.71826, 37.87939, 3.2159226, 0.037120353, -846.1443, 35.82311, 3.2159326, 0.041067485, -863.5399, 33.757996, 3.2128851, 0.044927154, -879.9012, 31.686125, 3.206821, 0.048696768, -895.2252, 29.609549, 3.1977825, 0.052373838, -909.51025, 27.530298, 3.1858149, 0.05595601, -922.75543, 25.450384, 3.1709654, 0.059441045, -934.9609, 23.371792, 3.1532838, 0.06282682, -946.12775, 21.296482, 3.1328213, 0.066111326, -956.25824, 19.226383, 3.1096315, 0.069292694, -965.35535, 17.163404, 3.0837703, 0.07236916, -973.42316, 15.109415, 3.0552945, 0.07533909, -980.46655, 13.066261, 3.0242636, 0.07820096, -986.4915, 11.03575, 2.9907384, 0.08095338, -991.5047, 9.019657, 2.9547813, 0.083595075, -995.51385, 7.0197234, 2.9164562, 0.0861249, -998.5274, 5.0376506, 2.8758287, 0.088541806, -1000.55475, 3.075104, 2.8329659, 0.090844885, -1001.606, 1.1337103, 2.7879357, 0.09303336, -1001.69226, -0.7849449, 2.7408075, 0.09510654, -1000.82513, -2.6793163, 2.691652, 0.09706387},
		'{-743.8243, 45.974236, 3.1845877, 0.020513162, -766.31213, 43.9743, 3.1971812, 0.024781875, -787.7957, 41.9571, 3.206581, 0.028974663, -808.2667, 39.924755, 3.2128172, 0.033088468, -827.71826, 37.87939, 3.2159226, 0.037120353, -846.1443, 35.82311, 3.2159326, 0.041067485, -863.5399, 33.757996, 3.2128851, 0.044927154, -879.9012, 31.686125, 3.206821, 0.048696768, -895.2252, 29.609549, 3.1977825, 0.052373838, -909.51025, 27.530298, 3.1858149, 0.05595601, -922.75543, 25.450384, 3.1709654, 0.059441045, -934.9609, 23.371792, 3.1532838, 0.06282682, -946.12775, 21.296482, 3.1328213, 0.066111326, -956.25824, 19.226383, 3.1096315, 0.069292694, -965.35535, 17.163404, 3.0837703, 0.07236916, -973.42316, 15.109415, 3.0552945, 0.07533909, -980.46655, 13.066261, 3.0242636, 0.07820096, -986.4915, 11.03575, 2.9907384, 0.08095338, -991.5047, 9.019657, 2.9547813, 0.083595075, -995.51385, 7.0197234, 2.9164562, 0.0861249, -998.5274, 5.0376506, 2.8758287, 0.088541806, -1000.55475, 3.075104, 2.8329659, 0.090844885, -1001.606, 1.1337103, 2.7879357, 0.09303336, -1001.69226, -0.7849449, 2.7408075, 0.09510654, -1000.82513, -2.6793163, 2.691652, 0.09706387},
		'{-741.83435, 45.861446, 3.1145601, 0.2656197, -764.2799, 43.927692, 3.0076368, 0.25940147, -785.7689, 42.035126, 2.9027734, 0.2532713, -806.32184, 40.183224, 2.7999477, 0.24722889, -825.95886, 38.371468, 2.699138, 0.24127385, -844.6999, 36.59935, 2.6003213, 0.23540583, -862.5647, 34.86634, 2.5034757, 0.22962445, -879.5727, 33.171936, 2.4085786, 0.22392929, -895.743, 31.515614, 2.3156075, 0.2183199, -911.09454, 29.89686, 2.2245402, 0.21279582, -925.646, 28.315166, 2.1353538, 0.20735663, -939.41583, 26.770018, 2.0480258, 0.2020018, -952.42206, 25.260904, 1.9625337, 0.19673084, -964.6826, 23.787321, 1.8788545, 0.1915432, -976.2152, 22.348759, 1.7969657, 0.18643838, -987.0372, 20.944714, 1.7168448, 0.18141583, -997.1656, 19.574684, 1.638469, 0.17647494, -1006.61743, 18.238169, 1.5618157, 0.17161517, -1015.40924, 16.934671, 1.4868623, 0.16683589, -1023.5575, 15.663694, 1.4135864, 0.16213652, -1031.0782, 14.424747, 1.3419652, 0.15751645, -1037.9875, 13.21734, 1.2719765, 0.15297502, -1044.3008, 12.040984, 1.2035977, 0.14851162, -1050.0336, 10.895195, 1.1368065, 0.14412557, -1055.201, 9.779492, 1.0715808, 0.13981622},
		'{-741.83435, 45.861446, 3.1145601, 0.2656197, -764.2799, 43.927692, 3.0076368, 0.25940147, -785.7689, 42.035126, 2.9027734, 0.2532713, -806.32184, 40.183224, 2.7999477, 0.24722889, -825.95886, 38.371468, 2.699138, 0.24127385, -844.6999, 36.59935, 2.6003213, 0.23540583, -862.5647, 34.86634, 2.5034757, 0.22962445, -879.5727, 33.171936, 2.4085786, 0.22392929, -895.743, 31.515614, 2.3156075, 0.2183199, -911.09454, 29.89686, 2.2245402, 0.21279582, -925.646, 28.315166, 2.1353538, 0.20735663, -939.41583, 26.770018, 2.0480258, 0.2020018, -952.42206, 25.260904, 1.9625337, 0.19673084, -964.6826, 23.787321, 1.8788545, 0.1915432, -976.2152, 22.348759, 1.7969657, 0.18643838, -987.0372, 20.944714, 1.7168448, 0.18141583, -997.1656, 19.574684, 1.638469, 0.17647494, -1006.61743, 18.238169, 1.5618157, 0.17161517, -1015.40924, 16.934671, 1.4868623, 0.16683589, -1023.5575, 15.663694, 1.4135864, 0.16213652, -1031.0782, 14.424747, 1.3419652, 0.15751645, -1037.9875, 13.21734, 1.2719765, 0.15297502, -1044.3008, 12.040984, 1.2035977, 0.14851162, -1050.0336, 10.895195, 1.1368065, 0.14412557, -1055.201, 9.779492, 1.0715808, 0.13981622}};
	localparam real Fbi[0:3][0:99] = '{
		'{909.9477, 56.318283, -1.1170552, -0.14624423, 881.5327, 57.330624, -1.0137653, -0.1446599, 852.62823, 58.276043, -0.91077894, -0.1429575, 823.2678, 59.154465, -0.8081901, -0.14114006, 793.4849, 59.965878, -0.70609146, -0.13921075, 763.3131, 60.710327, -0.6045741, -0.13717276, 732.78577, 61.387928, -0.5037274, -0.13502938, 701.9363, 61.99886, -0.40363896, -0.1327839, 670.798, 62.543354, -0.3043947, -0.13043976, 639.40393, 63.021717, -0.20607851, -0.12800038, 607.78723, 63.434296, -0.10877256, -0.12546922, 575.9805, 63.78151, -0.0125569245, -0.12284985, 544.01654, 64.06383, 0.0824903, -0.12014582, 511.92746, 64.281784, 0.1762931, -0.11736075, 479.74536, 64.43596, 0.26877755, -0.11449827, 447.502, 64.52698, 0.35987192, -0.111562066, 415.22882, 64.55554, 0.44950667, -0.108555816, 382.95676, 64.522385, 0.53761446, -0.10548326, 350.71658, 64.4283, 0.6241303, -0.102348104, 318.53848, 64.27412, 0.70899147, -0.09915412, 286.45233, 64.06072, 0.79213756, -0.09590506, 254.48747, 63.789047, 0.87351054, -0.09260468, 222.67284, 63.460064, 0.9530549, -0.089256756, 191.03679, 63.074787, 1.0307175, -0.08586505, 159.60725, 62.634277, 1.1064473, -0.08243332},
		'{-909.9477, -56.318283, 1.1170552, 0.14624423, -881.5327, -57.330624, 1.0137653, 0.1446599, -852.62823, -58.276043, 0.91077894, 0.1429575, -823.2678, -59.154465, 0.8081901, 0.14114006, -793.4849, -59.965878, 0.70609146, 0.13921075, -763.3131, -60.710327, 0.6045741, 0.13717276, -732.78577, -61.387928, 0.5037274, 0.13502938, -701.9363, -61.99886, 0.40363896, 0.1327839, -670.798, -62.543354, 0.3043947, 0.13043976, -639.40393, -63.021717, 0.20607851, 0.12800038, -607.78723, -63.434296, 0.10877256, 0.12546922, -575.9805, -63.78151, 0.0125569245, 0.12284985, -544.01654, -64.06383, -0.0824903, 0.12014582, -511.92746, -64.281784, -0.1762931, 0.11736075, -479.74536, -64.43596, -0.26877755, 0.11449827, -447.502, -64.52698, -0.35987192, 0.111562066, -415.22882, -64.55554, -0.44950667, 0.108555816, -382.95676, -64.522385, -0.53761446, 0.10548326, -350.71658, -64.4283, -0.6241303, 0.102348104, -318.53848, -64.27412, -0.70899147, 0.09915412, -286.45233, -64.06072, -0.79213756, 0.09590506, -254.48747, -63.789047, -0.87351054, 0.09260468, -222.67284, -63.460064, -0.9530549, 0.089256756, -191.03679, -63.074787, -1.0307175, 0.08586505, -159.60725, -62.634277, -1.1064473, 0.08243332},
		'{2770.766, 102.199974, 4.9312606, 0.18171343, 2719.9124, 101.213486, 4.894612, 0.1821949, 2669.554, 100.21841, 4.857218, 0.1825936, 2619.6953, 99.21537, 4.819115, 0.18291183, 2570.3398, 98.204994, 4.780339, 0.18315186, 2521.4915, 97.187874, 4.7409244, 0.18331595, 2473.153, 96.1646, 4.700905, 0.18340631, 2425.328, 95.13572, 4.6603136, 0.18342508, 2378.018, 94.10181, 4.619183, 0.1833744, 2331.2268, 93.0634, 4.577544, 0.18325639, 2284.9553, 92.02101, 4.5354285, 0.18307306, 2239.2063, 90.97515, 4.492866, 0.18282644, 2193.9807, 89.92633, 4.4498854, 0.18251851, 2149.2803, 88.875015, 4.4065156, 0.18215123, 2105.1062, 87.821686, 4.362785, 0.1817265, 2061.459, 86.76679, 4.31872, 0.18124618, 2018.3395, 85.710785, 4.274348, 0.18071212, 1975.7483, 84.654076, 4.2296934, 0.18012613, 1933.6854, 83.59711, 4.184783, 0.17948996, 1892.1511, 82.54026, 4.1396403, 0.17880537, 1851.1451, 81.48395, 4.0942893, 0.17807403, 1810.667, 80.428535, 4.0487537, 0.17729764, 1770.7163, 79.3744, 4.0030556, 0.17647782, 1731.2924, 78.3219, 3.9572175, 0.17561617, 1692.3942, 77.27138, 3.9112604, 0.17471428},
		'{-2770.766, -102.199974, -4.9312606, -0.18171343, -2719.9124, -101.213486, -4.894612, -0.1821949, -2669.554, -100.21841, -4.857218, -0.1825936, -2619.6953, -99.21537, -4.819115, -0.18291183, -2570.3398, -98.204994, -4.780339, -0.18315186, -2521.4915, -97.187874, -4.7409244, -0.18331595, -2473.153, -96.1646, -4.700905, -0.18340631, -2425.328, -95.13572, -4.6603136, -0.18342508, -2378.018, -94.10181, -4.619183, -0.1833744, -2331.2268, -93.0634, -4.577544, -0.18325639, -2284.9553, -92.02101, -4.5354285, -0.18307306, -2239.2063, -90.97515, -4.492866, -0.18282644, -2193.9807, -89.92633, -4.4498854, -0.18251851, -2149.2803, -88.875015, -4.4065156, -0.18215123, -2105.1062, -87.821686, -4.362785, -0.1817265, -2061.459, -86.76679, -4.31872, -0.18124618, -2018.3395, -85.710785, -4.274348, -0.18071212, -1975.7483, -84.654076, -4.2296934, -0.18012613, -1933.6854, -83.59711, -4.184783, -0.17948996, -1892.1511, -82.54026, -4.1396403, -0.17880537, -1851.1451, -81.48395, -4.0942893, -0.17807403, -1810.667, -80.428535, -4.0487537, -0.17729764, -1770.7163, -79.3744, -4.0030556, -0.17647782, -1731.2924, -78.3219, -3.9572175, -0.17561617, -1692.3942, -77.27138, -3.9112604, -0.17471428}};
	localparam real hf[0:1199] = {0.0104479985, -4.141178e-06, -5.3745443e-06, 4.2119637e-09, 0.010443858, -1.2420256e-05, -5.365872e-06, 1.2626676e-08, 0.01043558, -2.0689506e-05, -5.3485414e-06, 2.1014026e-08, 0.010423171, -2.894239e-05, -5.322578e-06, 2.9356382e-08, 0.010406641, -3.717239e-05, -5.288021e-06, 3.7636642e-08, 0.010386003, -4.537302e-05, -5.24492e-06, 4.5838235e-08, 0.010361274, -5.353783e-05, -5.1933366e-06, 5.3945122e-08, 0.010332473, -6.166041e-05, -5.133345e-06, 6.194182e-08, 0.010299622, -6.973439e-05, -5.0650283e-06, 6.981338e-08, 0.010262747, -7.775349e-05, -4.9884816e-06, 7.7545415e-08, 0.010221879, -8.571146e-05, -4.903811e-06, 8.512407e-08, 0.010177047, -9.360214e-05, -4.8111306e-06, 9.253608e-08, 0.0101282885, -0.00010141944, -4.710567e-06, 9.976869e-08, 0.010075641, -0.000109157365, -4.6022537e-06, 1.0680974e-07, 0.010019146, -0.00011681, -4.486335e-06, 1.13647616e-07, 0.0099588465, -0.00012437154, -4.362963e-06, 1.2027125e-07, 0.00989479, -0.00013183625, -4.2322995e-06, 1.2667016e-07, 0.009827027, -0.00013919856, -4.0945133e-06, 1.3283439e-07, 0.00975561, -0.00014645295, -3.949781e-06, 1.3875454e-07, 0.009680593, -0.00015359408, -3.7982875e-06, 1.4442182e-07, 0.009602035, -0.00016061669, -3.640224e-06, 1.4982791e-07, 0.009519997, -0.00016751567, -3.4757886e-06, 1.5496511e-07, 0.009434541, -0.00017428602, -3.3051863e-06, 1.598262e-07, 0.009345733, -0.00018092293, -3.128628e-06, 1.6440457e-07, 0.009253641, -0.00018742167, -2.9463297e-06, 1.686941e-07, 0.009158336, -0.00019377768, -2.7585136e-06, 1.7268921e-07, 0.009059888, -0.00019998659, -2.5654065e-06, 1.7638489e-07, 0.008958374, -0.00020604413, -2.3672399e-06, 1.7977658e-07, 0.0088538695, -0.00021194622, -2.16425e-06, 1.8286032e-07, 0.0087464545, -0.0002176889, -1.9566764e-06, 1.8563259e-07, 0.008636208, -0.00022326842, -1.7447629e-06, 1.8809043e-07, 0.008523214, -0.00022868118, -1.5287566e-06, 1.9023135e-07, 0.0084075555, -0.00023392374, -1.308907e-06, 1.9205335e-07, 0.0082893185, -0.00023899284, -1.085467e-06, 1.9355494e-07, 0.008168592, -0.0002438854, -8.586913e-07, 1.9473507e-07, 0.008045463, -0.0002485985, -6.2883686e-07, 1.9559319e-07, 0.007920024, -0.0002531294, -3.961621e-07, 1.9612919e-07, 0.007792365, -0.00025747553, -1.6092694e-07, 1.9634344e-07, 0.0076625794, -0.00026163453, 7.660774e-08, 1.962367e-07, 0.0075307614, -0.0002656042, 3.161804e-07, 1.9581022e-07, 0.0073970067, -0.00026938255, 5.5752906e-07, 1.9506562e-07, 0.0072614113, -0.00027296768, 8.0039166e-07, 1.9400498e-07, 0.007124072, -0.000276358, 1.0445063e-06, 1.9263078e-07, 0.006985086, -0.000279552, 1.289612e-06, 1.9094584e-07, 0.0068445527, -0.00028254843, 1.5354477e-06, 1.8895342e-07, 0.0067025707, -0.00028534618, 1.7817545e-06, 1.8665715e-07, 0.0065592397, -0.0002879443, 2.0282741e-06, 1.8406098e-07, 0.00641466, -0.00029034208, 2.2747502e-06, 1.8116924e-07, 0.006268931, -0.00029253896, 2.520928e-06, 1.7798662e-07, 0.006122154, -0.00029453455, 2.766556e-06, 1.7451808e-07, 0.00597443, -0.00029632865, 3.0113836e-06, 1.7076894e-07, 0.0058258595, -0.00029792127, 3.255164e-06, 1.6674484e-07, 0.0056765424, -0.00029931258, 3.497653e-06, 1.6245166e-07, 0.0055265804, -0.00030050287, 3.7386098e-06, 1.578956e-07, 0.005376073, -0.00030149266, 3.9777965e-06, 1.5308312e-07, 0.005225121, -0.00030228263, 4.214979e-06, 1.4802094e-07, 0.0050738235, -0.00030287364, 4.4499275e-06, 1.4271603e-07, 0.00492228, -0.0003032667, 4.6824152e-06, 1.3717559e-07, 0.0047705895, -0.00030346296, 4.9122214e-06, 1.3140702e-07, 0.0046188496, -0.0003034638, 5.1391285e-06, 1.2541798e-07, 0.004467158, -0.00030327073, 5.3629233e-06, 1.192163e-07, 0.004315611, -0.0003028854, 5.583398e-06, 1.1280996e-07, 0.0041643046, -0.0003023096, 5.8003498e-06, 1.06207175e-07, 0.004013333, -0.00030154534, 6.0135812e-06, 9.94163e-08, 0.0038627903, -0.00030059466, 6.2228996e-06, 9.2445816e-08, 0.003712769, -0.0002994599, 6.4281185e-06, 8.530438e-08, 0.0035633605, -0.00029814342, 6.6290563e-06, 7.800074e-08, 0.0034146553, -0.00029664775, 6.825537e-06, 7.054378e-08, 0.0032667422, -0.00029497556, 7.0173924e-06, 6.294247e-08, 0.0031197087, -0.00029312968, 7.2044572e-06, 5.5205888e-08, 0.002973641, -0.000291113, 7.3865745e-06, 4.734318e-08, 0.0028286236, -0.00028892866, 7.5635926e-06, 3.936356e-08, 0.00268474, -0.0002865797, 7.735367e-06, 3.1276297e-08, 0.0025420708, -0.00028406948, 7.901759e-06, 2.3090703e-08, 0.0024006967, -0.00028140142, 8.062636e-06, 1.481613e-08, 0.0022606952, -0.00027857895, 8.217873e-06, 6.4619448e-09, 0.0021221428, -0.00027560574, 8.36735e-06, -1.9624715e-09, 0.001985114, -0.00027248546, 8.510955e-06, -1.0447738e-08, 0.0018496813, -0.00026922193, 8.648583e-06, -1.8984483e-08, 0.0017159153, -0.000265819, 8.7801345e-06, -2.7563356e-08, 0.0015838848, -0.0002622807, 8.9055175e-06, -3.6175038e-08, 0.0014536565, -0.00025861102, 9.024647e-06, -4.481025e-08, 0.001325295, -0.00025481413, 9.137443e-06, -5.345976e-08, 0.0011988629, -0.00025089426, 9.243835e-06, -6.21144e-08, 0.0010744205, -0.0002468556, 9.343759e-06, -7.076508e-08, 0.00095202634, -0.00024270252, 9.437155e-06, -7.940278e-08, 0.00083173637, -0.00023843942, 9.523975e-06, -8.801856e-08, 0.0007136045, -0.00023407073, 9.604171e-06, -9.660358e-08, 0.0005976825, -0.00022960093, 9.6777085e-06, -1.0514913e-07, 0.0004840197, -0.00022503457, 9.7445545e-06, -1.1364657e-07, 0.00037266326, -0.00022037623, 9.804687e-06, -1.2208743e-07, 0.00026365803, -0.0002156305, 9.858087e-06, -1.3046333e-07, 0.00015704655, -0.00021080201, 9.904744e-06, -1.3876604e-07, 5.2869025e-05, -0.00020589546, 9.944654e-06, -1.4698749e-07, -4.883668e-05, -0.00020091551, 9.977821e-06, -1.5511975e-07, -0.00014803505, -0.00019586689, 1.0004252e-05, -1.6315502e-07, -0.0002446929, -0.00019075428, 1.0023962e-05, -1.7108573e-07, -0.00033877944, -0.00018558242, 1.0036973e-05, -1.789044e-07, -0.00043026623, -0.00018035604, 1.0043314e-05, -1.8660381e-07, -0.0005191272, -0.00017507988, 1.0043017e-05, -1.9417688e-07, -0.0006053386, -0.00016975864, 1.0036123e-05, -2.0161669e-07, -0.0006888791, -0.00016439703, 1.0022677e-05, -2.0891657e-07, -0.0007697297, -0.00015899977, 1.0002731e-05, -2.1607002e-07, -0.00084787374, -0.00015357153, 9.976342e-06, -2.2307077e-07, -0.00092329684, -0.00014811696, 9.943573e-06, -2.299127e-07, -0.0009959871, -0.0001426407, 9.904493e-06, -2.3658995e-07, -0.0010659347, -0.00013714736, 9.8591745e-06, -2.430969e-07, -0.0011331324, -0.0001316415, 9.807697e-06, -2.4942807e-07, -0.0011975749, -0.00012612766, 9.750145e-06, -2.5557827e-07, -0.0012592594, -0.000120610326, 9.686608e-06, -2.6154248e-07, -0.0013181854, -0.00011509395, 9.617179e-06, -2.67316e-07, -0.0013743542, -0.00010958292, 9.5419555e-06, -2.7289428e-07, -0.0014277699, -0.0001040816, 9.461043e-06, -2.78273e-07, -0.0014784381, -9.859427e-05, 9.3745475e-06, -2.8344814e-07, -0.0015263672, -9.3125156e-05, 9.282581e-06, -2.8841586e-07, -0.001571567, -8.767844e-05, 9.185259e-06, -2.9317258e-07, -0.00161405, -8.225823e-05, 9.0827025e-06, -2.9771496e-07, -0.0016538304, -7.686855e-05, 8.975034e-06, -3.020399e-07, -0.0016909243, -7.151338e-05, 8.86238e-06, -3.0614453e-07, -0.0017253502, -6.619661e-05, 8.7448725e-06, -3.1002625e-07, -0.0017571279, -6.0922055e-05, 8.6226455e-06, -3.1368268e-07, -0.0017862798, -5.5693454e-05, 8.4958365e-06, -3.1711167e-07, -0.0018128298, -5.051446e-05, 8.364584e-06, -3.2031136e-07, -0.0018368032, -4.5388653e-05, 8.229032e-06, -3.2328003e-07, -0.0018582278, -4.031951e-05, 8.089325e-06, -3.2601636e-07, -0.0018771327, -3.5310433e-05, 7.945613e-06, -3.285191e-07, -0.0018935488, -3.036473e-05, 7.798046e-06, -3.3078737e-07, -0.0019075086, -2.5485611e-05, 7.646774e-06, -3.328204e-07, -0.001919046, -2.0676196e-05, 7.491955e-06, -3.3461782e-07, -0.0019281969, -1.593951e-05, 7.3337433e-06, -3.361793e-07, -0.0019349981, -1.12784755e-05, 7.1722975e-06, -3.3750493e-07, -0.0019394885, -6.6959187e-06, 7.0077763e-06, -3.3859484e-07, -0.0019417076, -2.1945632e-06, 6.8403415e-06, -3.3944957e-07, -0.001941697, 2.2229692e-06, 6.6701546e-06, -3.4006973e-07, -0.001939499, 6.5541603e-06, 6.4973783e-06, -3.4045624e-07, -0.0019351576, 1.0796597e-05, 6.3221764e-06, -3.4061017e-07, -0.0019287176, 1.4947972e-05, 6.1447136e-06, -3.405329e-07, -0.0019202251, 1.9006084e-05, 5.9651543e-06, -3.4022594e-07, -0.0019097273, 2.296884e-05, 5.7836633e-06, -3.3969098e-07, -0.0018972725, 2.6834254e-05, 5.600407e-06, -3.3893002e-07, -0.0018829097, 3.060045e-05, 5.41555e-06, -3.3794518e-07, -0.001866689, 3.4265664e-05, 5.229257e-06, -3.367388e-07, -0.0018486611, 3.782823e-05, 5.0416943e-06, -3.3531336e-07, -0.0018288781, 4.128661e-05, 4.853025e-06, -3.3367158e-07, -0.0018073921, 4.463936e-05, 4.663414e-06, -3.3181635e-07, -0.0017842565, 4.7885154e-05, 4.473023e-06, -3.2975075e-07, -0.001759525, 5.1022773e-05, 4.2820157e-06, -3.2747798e-07, -0.001733252, 5.405111e-05, 4.090552e-06, -3.2500148e-07, -0.0017054923, 5.6969166e-05, 3.8987923e-06, -3.2232475e-07, -0.0016763014, 5.977605e-05, 3.7068953e-06, -3.1945157e-07, -0.0016457349, 6.247099e-05, 3.515018e-06, -3.1638575e-07, -0.0016138491, 6.50533e-05, 3.3233162e-06, -3.1313132e-07, -0.0015807004, 6.7522415e-05, 3.1319432e-06, -3.0969244e-07, -0.0015463457, 6.987788e-05, 2.9410517e-06, -3.060734e-07, -0.0015108415, 7.211936e-05, 2.750791e-06, -3.0227858e-07, -0.0014742453, 7.424658e-05, 2.5613097e-06, -2.9831256e-07, -0.0014366141, 7.625941e-05, 2.3727532e-06, -2.9417996e-07, -0.0013980049, 7.815781e-05, 2.185265e-06, -2.8988555e-07, -0.0013584753, 7.994185e-05, 1.998986e-06, -2.8543423e-07, -0.0013180822, 8.1611666e-05, 1.8140547e-06, -2.8083096e-07, -0.0012768826, 8.316754e-05, 1.6306071e-06, -2.7608078e-07, -0.0012349335, 8.460983e-05, 1.4487763e-06, -2.711889e-07, -0.0011922916, 8.593898e-05, 1.2686925e-06, -2.661605e-07, -0.0011490133, 8.7155546e-05, 1.090483e-06, -2.610009e-07, -0.0011051547, 8.8260174e-05, 9.142722e-07, -2.5571555e-07, -0.0010607716, 8.925359e-05, 7.401815e-07, -2.5030985e-07, -0.0010159196, 9.013662e-05, 5.683289e-07, -2.4478933e-07, -0.0009706533, 9.091018e-05, 3.988293e-07, -2.3915953e-07, -0.0009250275, 9.157527e-05, 2.317942e-07, -2.3342606e-07, -0.0008790959, 9.213296e-05, 6.733187e-08, -2.2759461e-07, -0.0008329122, 9.258442e-05, -9.445301e-08, -2.2167083e-07, -0.00078652904, 9.2930895e-05, -2.534592e-07, -2.1566046e-07, -0.0007399986, 9.317371e-05, -4.0958903e-07, -2.0956922e-07, -0.0006933724, 9.3314244e-05, -5.627485e-07, -2.034029e-07, -0.00064670114, 9.3353985e-05, -7.1284705e-07, -1.9716725e-07, -0.00060003495, 9.329447e-05, -8.5979815e-07, -1.9086805e-07, -0.00055342296, 9.313731e-05, -1.0035188e-06, -1.845111e-07, -0.00050691364, 9.288418e-05, -1.1439298e-06, -1.7810216e-07, -0.00046055447, 9.2536815e-05, -1.2809558e-06, -1.7164699e-07, -0.0004143922, 9.209703e-05, -1.4145252e-06, -1.6515136e-07, -0.00036847254, 9.156668e-05, -1.5445704e-06, -1.58621e-07, -0.0003228403, 9.0947695e-05, -1.6710276e-06, -1.5206162e-07, -0.0002775393, 9.0242036e-05, -1.7938369e-06, -1.454789e-07, -0.00023261236, 8.945174e-05, -1.9129423e-06, -1.3887846e-07, -0.00018810132, 8.857889e-05, -2.0282916e-06, -1.3226592e-07, -0.00014404689, 8.7625594e-05, -2.1398369e-06, -1.2564684e-07, -0.00010048877, 8.659403e-05, -2.2475338e-06, -1.1902671e-07, -5.7465535e-05, 8.5486405e-05, -2.351342e-06, -1.1241099e-07, -1.5014663e-05, 8.430497e-05, -2.451225e-06, -1.0580507e-07, 2.6827514e-05, 8.3052015e-05, -2.5471506e-06, -9.921428e-08, 6.8025816e-05, 8.172986e-05, -2.6390899e-06, -9.264389e-08, 0.00010854623, 8.034085e-05, -2.727018e-06, -8.609907e-08, 0.00014835592, 7.888738e-05, -2.8109143e-06, -7.958494e-08, 0.00018742327, 7.737186e-05, -2.8907618e-06, -7.3106534e-08, 0.00022571784, 7.579671e-05, -2.9665468e-06, -6.6668804e-08, 0.00026321044, 7.416439e-05, -3.03826e-06, -6.02766e-08, 0.00029987312, 7.2477385e-05, -3.1058958e-06, -5.393469e-08, 0.00033567913, 7.073818e-05, -3.169452e-06, -4.7647756e-08, 0.000370603, 6.894927e-05, -3.2289297e-06, -4.1420368e-08, 0.00040462054, 6.711319e-05, -3.2843345e-06, -3.5257003e-08, 0.00043770878, 6.523246e-05, -3.3356753e-06, -2.9162026e-08, 0.00046984598, 6.3309606e-05, -3.3829638e-06, -2.3139702e-08, 0.0005010118, 6.134717e-05, -3.4262162e-06, -1.7194179e-08, 0.000531187, 5.9347687e-05, -3.465451e-06, -1.1329499e-08, 0.0005603537, 5.73137e-05, -3.5006915e-06, -5.5495843e-09, 0.00058849534, 5.5247743e-05, -3.5319626e-06, 1.4176046e-10, 0.00061559654, 5.3152344e-05, -3.559294e-06, 5.7408505e-09, 0.0006416432, 5.1030027e-05, -3.5827175e-06, 1.1244122e-08, 0.0006666225, 4.888331e-05, -3.6022682e-06, 1.6648137e-08, 0.00069052284, 4.671469e-05, -3.6179847e-06, 2.1949583e-08, 0.00071333395, 4.4526656e-05, -3.629908e-06, 2.7145276e-08, 0.0007350467, 4.2321677e-05, -3.6380823e-06, 3.223216e-08, 0.0007556532, 4.010221e-05, -3.6425545e-06, 3.7207304e-08, 0.0007751469, 3.7870686e-05, -3.6433744e-06, 4.2067924e-08, 0.0007935223, 3.5629517e-05, -3.6405943e-06, 4.681136e-08, 0.0008107752, 3.3381086e-05, -3.634269e-06, 5.1435077e-08, 0.0008269026, 3.1127754e-05, -3.624456e-06, 5.5936688e-08, 0.0008419025, 2.8871857e-05, -3.6112153e-06, 6.0313944e-08, 0.0008557744, 2.6615695e-05, -3.5946086e-06, 6.4564716e-08, 0.00086851855, 2.4361538e-05, -3.574701e-06, 6.868703e-08, 0.0008801366, 2.2111624e-05, -3.5515584e-06, 7.2679036e-08, 0.0008906312, 1.9868156e-05, -3.5252497e-06, 7.6539024e-08, 0.0009000062, 1.76333e-05, -3.4958457e-06, 8.026543e-08, 0.00090826635, 1.5409183e-05, -3.4634188e-06, 8.385681e-08, 0.0009154175, 1.3197895e-05, -3.4280433e-06, 8.7311875e-08, 0.00092146674, 1.1001483e-05, -3.3897954e-06, 9.0629456e-08, 0.00092642184, 8.82195e-06, -3.3487527e-06, 9.380853e-08, 0.0009302918, 6.66126e-06, -3.3049944e-06, 9.684821e-08, 0.00093308656, 4.521327e-06, -3.258601e-06, 9.9747744e-08, 0.0009348169, 2.4040214e-06, -3.2096552e-06, 1.0250651e-07, 0.00093549467, 3.1116593e-07, -3.1582395e-06, 1.05124016e-07, 0.00093513244, -1.7554657e-06, -3.104439e-06, 1.075999e-07, 0.00093374384, -3.794149e-06, -3.0483386e-06, 1.0993395e-07, 0.00093134324, -5.8032097e-06, -2.9900255e-06, 1.1212607e-07, 0.00092794583, -7.7810255e-06, -2.9295866e-06, 1.14176274e-07, 0.0009235677, -9.726027e-06, -2.8671104e-06, 1.16084735e-07, 0.0009182255, -1.16366955e-05, -2.802686e-06, 1.1785174e-07, 0.0009119369, -1.3511569e-05, -2.7364024e-06, 1.1947768e-07, 0.00090472016, -1.5349236e-05, -2.6683504e-06, 1.209631e-07, 0.00089659414, -1.7148348e-05, -2.5986199e-06, 1.2230863e-07, 0.00088757847, -1.8907602e-05, -2.527302e-06, 1.2351505e-07, 0.00087769335, -2.0625757e-05, -2.4544881e-06, 1.2458324e-07, 0.00086695974, -2.230163e-05, -2.3802693e-06, 1.2551418e-07, 0.000855399, -2.3934092e-05, -2.3047369e-06, 1.2630899e-07, 0.0008430331, -2.552207e-05, -2.2279826e-06, 1.2696887e-07, 0.0008298845, -2.7064552e-05, -2.1500975e-06, 1.2749514e-07, 0.00081597624, -2.8560584e-05, -2.071173e-06, 1.2788924e-07, 0.00080133183, -3.0009267e-05, -1.9913e-06, 1.2815268e-07, 0.000785975, -3.1409763e-05, -1.910569e-06, 1.282871e-07, 0.0007699302, -3.2761287e-05, -1.8290699e-06, 1.2829419e-07, 0.00075322203, -3.406312e-05, -1.746893e-06, 1.281758e-07, 0.00073587545, -3.531459e-05, -1.6641271e-06, 1.2793382e-07, 0.00071791594, -3.6515103e-05, -1.5808608e-06, 1.2757022e-07, 0.00069936895, -3.7664096e-05, -1.497182e-06, 1.270871e-07, 0.0006802605, -3.876108e-05, -1.4131775e-06, 1.2648664e-07, 0.0006606166, -3.9805625e-05, -1.3289335e-06, 1.2577102e-07, 0.00064046367, -4.079735e-05, -1.2445354e-06, 1.2494262e-07, 0.0006198281, -4.1735933e-05, -1.1600672e-06, 1.2400376e-07, 0.00059873663, -4.2621108e-05, -1.0756123e-06, 1.2295696e-07, 0.000577216, -4.3452666e-05, -9.912526e-07, 1.218047e-07, 0.00055529294, -4.4230455e-05, -9.070691e-07, 1.2054959e-07, 0.00053299445, -4.495437e-05, -8.231413e-07, 1.1919426e-07, 0.00051034754, -4.562437e-05, -7.3954754e-07, 1.1774143e-07, 0.0004873791, -4.6240453e-05, -6.563648e-07, 1.1619386e-07, 0.00046411608, -4.680269e-05, -5.7366873e-07, 1.14554354e-07, 0.00044058537, -4.7311183e-05, -4.915332e-07, 1.12825774e-07, 0.00041681383, -4.77661e-05, -4.100309e-07, 1.11011026e-07, 0.00039282817, -4.816765e-05, -3.292328e-07, 1.09113046e-07, 0.00036865502, -4.85161e-05, -2.4920823e-07, 1.07134824e-07, 0.00034432087, -4.8811755e-05, -1.7002498e-07, 1.0507937e-07, 0.000319852, -4.9054976e-05, -9.1749e-08, 1.0294975e-07, 0.00029527457, -4.924617e-05, -1.4444599e-08, 1.0074902e-07, 0.00027061443, -4.938578e-05, 6.182573e-08, 9.848029e-08, 0.0002458973, -4.9474307e-05, 1.3700131e-07, 9.61467e-08, 0.00022114856, -4.9512284e-05, 2.1102329e-07, 9.3751375e-08, 0.00019639333, -4.95003e-05, 2.8383474e-07, 9.129749e-08, 0.00017165647, -4.943897e-05, 3.5538062e-07, 8.8788205e-08, 0.00014696248, -4.9328963e-05, 4.256078e-07, 8.6226706e-08, 0.0001223355, -4.9170976e-05, 4.9446516e-07, 8.3616186e-08, 9.779938e-05, -4.8965747e-05, 5.619035e-07, 8.0959836e-08, 7.337751e-05, -4.8714057e-05, 6.278757e-07, 7.8260854e-08, 4.909293e-05, -4.8416714e-05, 6.923366e-07, 7.552242e-08, 2.496826e-05, -4.807457e-05, 7.5524315e-07, 7.2747724e-08, 1.0256822e-06, -4.7688496e-05, 8.1655435e-07, 6.9939944e-08, -2.2713066e-05, -4.7259407e-05, 8.762311e-07, 6.710225e-08, -4.6226713e-05, -4.6788246e-05, 9.342367e-07, 6.423778e-08, -6.949446e-05, -4.627598e-05, 9.905363e-07, 6.134968e-08, -9.249601e-05, -4.5723613e-05, 1.0450971e-06, 5.844107e-08, -0.00011521156, -4.5132165e-05, 1.0978886e-06, 5.5515038e-08, -0.00013762184, -4.4502685e-05, 1.1488822e-06, 5.2574652e-08, -0.00015970808, -4.383625e-05, 1.1980516e-06, 4.9622958e-08, -0.00018145211, -4.3133958e-05, 1.2453723e-06, 4.666296e-08, -0.00020283625, -4.239692e-05, 1.2908224e-06, 4.3697653e-08, -0.00022384342, -4.1626285e-05, 1.3343815e-06, 4.0729972e-08, -0.00024445713, -4.08232e-05, 1.3760317e-06, 3.7762828e-08, -0.00026466142, -3.998884e-05, 1.415757e-06, 3.479909e-08, -0.00028444096, -3.9124403e-05, 1.4535434e-06, 3.184159e-08, -0.000303781, -3.823108e-05, 1.4893791e-06, 2.8893115e-08, -0.00032266742, -3.7310096e-05, 1.5232544e-06, 2.5956403e-08, -0.0003410867, -3.636268e-05, 1.5551611e-06, 2.3034145e-08};
	localparam real hb[0:1199] = {0.0104479985, 4.141178e-06, -5.3745443e-06, -4.2119637e-09, 0.010443858, 1.2420256e-05, -5.365872e-06, -1.2626676e-08, 0.01043558, 2.0689506e-05, -5.3485414e-06, -2.1014026e-08, 0.010423171, 2.894239e-05, -5.322578e-06, -2.9356382e-08, 0.010406641, 3.717239e-05, -5.288021e-06, -3.7636642e-08, 0.010386003, 4.537302e-05, -5.24492e-06, -4.5838235e-08, 0.010361274, 5.353783e-05, -5.1933366e-06, -5.3945122e-08, 0.010332473, 6.166041e-05, -5.133345e-06, -6.194182e-08, 0.010299622, 6.973439e-05, -5.0650283e-06, -6.981338e-08, 0.010262747, 7.775349e-05, -4.9884816e-06, -7.7545415e-08, 0.010221879, 8.571146e-05, -4.903811e-06, -8.512407e-08, 0.010177047, 9.360214e-05, -4.8111306e-06, -9.253608e-08, 0.0101282885, 0.00010141944, -4.710567e-06, -9.976869e-08, 0.010075641, 0.000109157365, -4.6022537e-06, -1.0680974e-07, 0.010019146, 0.00011681, -4.486335e-06, -1.13647616e-07, 0.0099588465, 0.00012437154, -4.362963e-06, -1.2027125e-07, 0.00989479, 0.00013183625, -4.2322995e-06, -1.2667016e-07, 0.009827027, 0.00013919856, -4.0945133e-06, -1.3283439e-07, 0.00975561, 0.00014645295, -3.949781e-06, -1.3875454e-07, 0.009680593, 0.00015359408, -3.7982875e-06, -1.4442182e-07, 0.009602035, 0.00016061669, -3.640224e-06, -1.4982791e-07, 0.009519997, 0.00016751567, -3.4757886e-06, -1.5496511e-07, 0.009434541, 0.00017428602, -3.3051863e-06, -1.598262e-07, 0.009345733, 0.00018092293, -3.128628e-06, -1.6440457e-07, 0.009253641, 0.00018742167, -2.9463297e-06, -1.686941e-07, 0.009158336, 0.00019377768, -2.7585136e-06, -1.7268921e-07, 0.009059888, 0.00019998659, -2.5654065e-06, -1.7638489e-07, 0.008958374, 0.00020604413, -2.3672399e-06, -1.7977658e-07, 0.0088538695, 0.00021194622, -2.16425e-06, -1.8286032e-07, 0.0087464545, 0.0002176889, -1.9566764e-06, -1.8563259e-07, 0.008636208, 0.00022326842, -1.7447629e-06, -1.8809043e-07, 0.008523214, 0.00022868118, -1.5287566e-06, -1.9023135e-07, 0.0084075555, 0.00023392374, -1.308907e-06, -1.9205335e-07, 0.0082893185, 0.00023899284, -1.085467e-06, -1.9355494e-07, 0.008168592, 0.0002438854, -8.586913e-07, -1.9473507e-07, 0.008045463, 0.0002485985, -6.2883686e-07, -1.9559319e-07, 0.007920024, 0.0002531294, -3.961621e-07, -1.9612919e-07, 0.007792365, 0.00025747553, -1.6092694e-07, -1.9634344e-07, 0.0076625794, 0.00026163453, 7.660774e-08, -1.962367e-07, 0.0075307614, 0.0002656042, 3.161804e-07, -1.9581022e-07, 0.0073970067, 0.00026938255, 5.5752906e-07, -1.9506562e-07, 0.0072614113, 0.00027296768, 8.0039166e-07, -1.9400498e-07, 0.007124072, 0.000276358, 1.0445063e-06, -1.9263078e-07, 0.006985086, 0.000279552, 1.289612e-06, -1.9094584e-07, 0.0068445527, 0.00028254843, 1.5354477e-06, -1.8895342e-07, 0.0067025707, 0.00028534618, 1.7817545e-06, -1.8665715e-07, 0.0065592397, 0.0002879443, 2.0282741e-06, -1.8406098e-07, 0.00641466, 0.00029034208, 2.2747502e-06, -1.8116924e-07, 0.006268931, 0.00029253896, 2.520928e-06, -1.7798662e-07, 0.006122154, 0.00029453455, 2.766556e-06, -1.7451808e-07, 0.00597443, 0.00029632865, 3.0113836e-06, -1.7076894e-07, 0.0058258595, 0.00029792127, 3.255164e-06, -1.6674484e-07, 0.0056765424, 0.00029931258, 3.497653e-06, -1.6245166e-07, 0.0055265804, 0.00030050287, 3.7386098e-06, -1.578956e-07, 0.005376073, 0.00030149266, 3.9777965e-06, -1.5308312e-07, 0.005225121, 0.00030228263, 4.214979e-06, -1.4802094e-07, 0.0050738235, 0.00030287364, 4.4499275e-06, -1.4271603e-07, 0.00492228, 0.0003032667, 4.6824152e-06, -1.3717559e-07, 0.0047705895, 0.00030346296, 4.9122214e-06, -1.3140702e-07, 0.0046188496, 0.0003034638, 5.1391285e-06, -1.2541798e-07, 0.004467158, 0.00030327073, 5.3629233e-06, -1.192163e-07, 0.004315611, 0.0003028854, 5.583398e-06, -1.1280996e-07, 0.0041643046, 0.0003023096, 5.8003498e-06, -1.06207175e-07, 0.004013333, 0.00030154534, 6.0135812e-06, -9.94163e-08, 0.0038627903, 0.00030059466, 6.2228996e-06, -9.2445816e-08, 0.003712769, 0.0002994599, 6.4281185e-06, -8.530438e-08, 0.0035633605, 0.00029814342, 6.6290563e-06, -7.800074e-08, 0.0034146553, 0.00029664775, 6.825537e-06, -7.054378e-08, 0.0032667422, 0.00029497556, 7.0173924e-06, -6.294247e-08, 0.0031197087, 0.00029312968, 7.2044572e-06, -5.5205888e-08, 0.002973641, 0.000291113, 7.3865745e-06, -4.734318e-08, 0.0028286236, 0.00028892866, 7.5635926e-06, -3.936356e-08, 0.00268474, 0.0002865797, 7.735367e-06, -3.1276297e-08, 0.0025420708, 0.00028406948, 7.901759e-06, -2.3090703e-08, 0.0024006967, 0.00028140142, 8.062636e-06, -1.481613e-08, 0.0022606952, 0.00027857895, 8.217873e-06, -6.4619448e-09, 0.0021221428, 0.00027560574, 8.36735e-06, 1.9624715e-09, 0.001985114, 0.00027248546, 8.510955e-06, 1.0447738e-08, 0.0018496813, 0.00026922193, 8.648583e-06, 1.8984483e-08, 0.0017159153, 0.000265819, 8.7801345e-06, 2.7563356e-08, 0.0015838848, 0.0002622807, 8.9055175e-06, 3.6175038e-08, 0.0014536565, 0.00025861102, 9.024647e-06, 4.481025e-08, 0.001325295, 0.00025481413, 9.137443e-06, 5.345976e-08, 0.0011988629, 0.00025089426, 9.243835e-06, 6.21144e-08, 0.0010744205, 0.0002468556, 9.343759e-06, 7.076508e-08, 0.00095202634, 0.00024270252, 9.437155e-06, 7.940278e-08, 0.00083173637, 0.00023843942, 9.523975e-06, 8.801856e-08, 0.0007136045, 0.00023407073, 9.604171e-06, 9.660358e-08, 0.0005976825, 0.00022960093, 9.6777085e-06, 1.0514913e-07, 0.0004840197, 0.00022503457, 9.7445545e-06, 1.1364657e-07, 0.00037266326, 0.00022037623, 9.804687e-06, 1.2208743e-07, 0.00026365803, 0.0002156305, 9.858087e-06, 1.3046333e-07, 0.00015704655, 0.00021080201, 9.904744e-06, 1.3876604e-07, 5.2869025e-05, 0.00020589546, 9.944654e-06, 1.4698749e-07, -4.883668e-05, 0.00020091551, 9.977821e-06, 1.5511975e-07, -0.00014803505, 0.00019586689, 1.0004252e-05, 1.6315502e-07, -0.0002446929, 0.00019075428, 1.0023962e-05, 1.7108573e-07, -0.00033877944, 0.00018558242, 1.0036973e-05, 1.789044e-07, -0.00043026623, 0.00018035604, 1.0043314e-05, 1.8660381e-07, -0.0005191272, 0.00017507988, 1.0043017e-05, 1.9417688e-07, -0.0006053386, 0.00016975864, 1.0036123e-05, 2.0161669e-07, -0.0006888791, 0.00016439703, 1.0022677e-05, 2.0891657e-07, -0.0007697297, 0.00015899977, 1.0002731e-05, 2.1607002e-07, -0.00084787374, 0.00015357153, 9.976342e-06, 2.2307077e-07, -0.00092329684, 0.00014811696, 9.943573e-06, 2.299127e-07, -0.0009959871, 0.0001426407, 9.904493e-06, 2.3658995e-07, -0.0010659347, 0.00013714736, 9.8591745e-06, 2.430969e-07, -0.0011331324, 0.0001316415, 9.807697e-06, 2.4942807e-07, -0.0011975749, 0.00012612766, 9.750145e-06, 2.5557827e-07, -0.0012592594, 0.000120610326, 9.686608e-06, 2.6154248e-07, -0.0013181854, 0.00011509395, 9.617179e-06, 2.67316e-07, -0.0013743542, 0.00010958292, 9.5419555e-06, 2.7289428e-07, -0.0014277699, 0.0001040816, 9.461043e-06, 2.78273e-07, -0.0014784381, 9.859427e-05, 9.3745475e-06, 2.8344814e-07, -0.0015263672, 9.3125156e-05, 9.282581e-06, 2.8841586e-07, -0.001571567, 8.767844e-05, 9.185259e-06, 2.9317258e-07, -0.00161405, 8.225823e-05, 9.0827025e-06, 2.9771496e-07, -0.0016538304, 7.686855e-05, 8.975034e-06, 3.020399e-07, -0.0016909243, 7.151338e-05, 8.86238e-06, 3.0614453e-07, -0.0017253502, 6.619661e-05, 8.7448725e-06, 3.1002625e-07, -0.0017571279, 6.0922055e-05, 8.6226455e-06, 3.1368268e-07, -0.0017862798, 5.5693454e-05, 8.4958365e-06, 3.1711167e-07, -0.0018128298, 5.051446e-05, 8.364584e-06, 3.2031136e-07, -0.0018368032, 4.5388653e-05, 8.229032e-06, 3.2328003e-07, -0.0018582278, 4.031951e-05, 8.089325e-06, 3.2601636e-07, -0.0018771327, 3.5310433e-05, 7.945613e-06, 3.285191e-07, -0.0018935488, 3.036473e-05, 7.798046e-06, 3.3078737e-07, -0.0019075086, 2.5485611e-05, 7.646774e-06, 3.328204e-07, -0.001919046, 2.0676196e-05, 7.491955e-06, 3.3461782e-07, -0.0019281969, 1.593951e-05, 7.3337433e-06, 3.361793e-07, -0.0019349981, 1.12784755e-05, 7.1722975e-06, 3.3750493e-07, -0.0019394885, 6.6959187e-06, 7.0077763e-06, 3.3859484e-07, -0.0019417076, 2.1945632e-06, 6.8403415e-06, 3.3944957e-07, -0.001941697, -2.2229692e-06, 6.6701546e-06, 3.4006973e-07, -0.001939499, -6.5541603e-06, 6.4973783e-06, 3.4045624e-07, -0.0019351576, -1.0796597e-05, 6.3221764e-06, 3.4061017e-07, -0.0019287176, -1.4947972e-05, 6.1447136e-06, 3.405329e-07, -0.0019202251, -1.9006084e-05, 5.9651543e-06, 3.4022594e-07, -0.0019097273, -2.296884e-05, 5.7836633e-06, 3.3969098e-07, -0.0018972725, -2.6834254e-05, 5.600407e-06, 3.3893002e-07, -0.0018829097, -3.060045e-05, 5.41555e-06, 3.3794518e-07, -0.001866689, -3.4265664e-05, 5.229257e-06, 3.367388e-07, -0.0018486611, -3.782823e-05, 5.0416943e-06, 3.3531336e-07, -0.0018288781, -4.128661e-05, 4.853025e-06, 3.3367158e-07, -0.0018073921, -4.463936e-05, 4.663414e-06, 3.3181635e-07, -0.0017842565, -4.7885154e-05, 4.473023e-06, 3.2975075e-07, -0.001759525, -5.1022773e-05, 4.2820157e-06, 3.2747798e-07, -0.001733252, -5.405111e-05, 4.090552e-06, 3.2500148e-07, -0.0017054923, -5.6969166e-05, 3.8987923e-06, 3.2232475e-07, -0.0016763014, -5.977605e-05, 3.7068953e-06, 3.1945157e-07, -0.0016457349, -6.247099e-05, 3.515018e-06, 3.1638575e-07, -0.0016138491, -6.50533e-05, 3.3233162e-06, 3.1313132e-07, -0.0015807004, -6.7522415e-05, 3.1319432e-06, 3.0969244e-07, -0.0015463457, -6.987788e-05, 2.9410517e-06, 3.060734e-07, -0.0015108415, -7.211936e-05, 2.750791e-06, 3.0227858e-07, -0.0014742453, -7.424658e-05, 2.5613097e-06, 2.9831256e-07, -0.0014366141, -7.625941e-05, 2.3727532e-06, 2.9417996e-07, -0.0013980049, -7.815781e-05, 2.185265e-06, 2.8988555e-07, -0.0013584753, -7.994185e-05, 1.998986e-06, 2.8543423e-07, -0.0013180822, -8.1611666e-05, 1.8140547e-06, 2.8083096e-07, -0.0012768826, -8.316754e-05, 1.6306071e-06, 2.7608078e-07, -0.0012349335, -8.460983e-05, 1.4487763e-06, 2.711889e-07, -0.0011922916, -8.593898e-05, 1.2686925e-06, 2.661605e-07, -0.0011490133, -8.7155546e-05, 1.090483e-06, 2.610009e-07, -0.0011051547, -8.8260174e-05, 9.142722e-07, 2.5571555e-07, -0.0010607716, -8.925359e-05, 7.401815e-07, 2.5030985e-07, -0.0010159196, -9.013662e-05, 5.683289e-07, 2.4478933e-07, -0.0009706533, -9.091018e-05, 3.988293e-07, 2.3915953e-07, -0.0009250275, -9.157527e-05, 2.317942e-07, 2.3342606e-07, -0.0008790959, -9.213296e-05, 6.733187e-08, 2.2759461e-07, -0.0008329122, -9.258442e-05, -9.445301e-08, 2.2167083e-07, -0.00078652904, -9.2930895e-05, -2.534592e-07, 2.1566046e-07, -0.0007399986, -9.317371e-05, -4.0958903e-07, 2.0956922e-07, -0.0006933724, -9.3314244e-05, -5.627485e-07, 2.034029e-07, -0.00064670114, -9.3353985e-05, -7.1284705e-07, 1.9716725e-07, -0.00060003495, -9.329447e-05, -8.5979815e-07, 1.9086805e-07, -0.00055342296, -9.313731e-05, -1.0035188e-06, 1.845111e-07, -0.00050691364, -9.288418e-05, -1.1439298e-06, 1.7810216e-07, -0.00046055447, -9.2536815e-05, -1.2809558e-06, 1.7164699e-07, -0.0004143922, -9.209703e-05, -1.4145252e-06, 1.6515136e-07, -0.00036847254, -9.156668e-05, -1.5445704e-06, 1.58621e-07, -0.0003228403, -9.0947695e-05, -1.6710276e-06, 1.5206162e-07, -0.0002775393, -9.0242036e-05, -1.7938369e-06, 1.454789e-07, -0.00023261236, -8.945174e-05, -1.9129423e-06, 1.3887846e-07, -0.00018810132, -8.857889e-05, -2.0282916e-06, 1.3226592e-07, -0.00014404689, -8.7625594e-05, -2.1398369e-06, 1.2564684e-07, -0.00010048877, -8.659403e-05, -2.2475338e-06, 1.1902671e-07, -5.7465535e-05, -8.5486405e-05, -2.351342e-06, 1.1241099e-07, -1.5014663e-05, -8.430497e-05, -2.451225e-06, 1.0580507e-07, 2.6827514e-05, -8.3052015e-05, -2.5471506e-06, 9.921428e-08, 6.8025816e-05, -8.172986e-05, -2.6390899e-06, 9.264389e-08, 0.00010854623, -8.034085e-05, -2.727018e-06, 8.609907e-08, 0.00014835592, -7.888738e-05, -2.8109143e-06, 7.958494e-08, 0.00018742327, -7.737186e-05, -2.8907618e-06, 7.3106534e-08, 0.00022571784, -7.579671e-05, -2.9665468e-06, 6.6668804e-08, 0.00026321044, -7.416439e-05, -3.03826e-06, 6.02766e-08, 0.00029987312, -7.2477385e-05, -3.1058958e-06, 5.393469e-08, 0.00033567913, -7.073818e-05, -3.169452e-06, 4.7647756e-08, 0.000370603, -6.894927e-05, -3.2289297e-06, 4.1420368e-08, 0.00040462054, -6.711319e-05, -3.2843345e-06, 3.5257003e-08, 0.00043770878, -6.523246e-05, -3.3356753e-06, 2.9162026e-08, 0.00046984598, -6.3309606e-05, -3.3829638e-06, 2.3139702e-08, 0.0005010118, -6.134717e-05, -3.4262162e-06, 1.7194179e-08, 0.000531187, -5.9347687e-05, -3.465451e-06, 1.1329499e-08, 0.0005603537, -5.73137e-05, -3.5006915e-06, 5.5495843e-09, 0.00058849534, -5.5247743e-05, -3.5319626e-06, -1.4176046e-10, 0.00061559654, -5.3152344e-05, -3.559294e-06, -5.7408505e-09, 0.0006416432, -5.1030027e-05, -3.5827175e-06, -1.1244122e-08, 0.0006666225, -4.888331e-05, -3.6022682e-06, -1.6648137e-08, 0.00069052284, -4.671469e-05, -3.6179847e-06, -2.1949583e-08, 0.00071333395, -4.4526656e-05, -3.629908e-06, -2.7145276e-08, 0.0007350467, -4.2321677e-05, -3.6380823e-06, -3.223216e-08, 0.0007556532, -4.010221e-05, -3.6425545e-06, -3.7207304e-08, 0.0007751469, -3.7870686e-05, -3.6433744e-06, -4.2067924e-08, 0.0007935223, -3.5629517e-05, -3.6405943e-06, -4.681136e-08, 0.0008107752, -3.3381086e-05, -3.634269e-06, -5.1435077e-08, 0.0008269026, -3.1127754e-05, -3.624456e-06, -5.5936688e-08, 0.0008419025, -2.8871857e-05, -3.6112153e-06, -6.0313944e-08, 0.0008557744, -2.6615695e-05, -3.5946086e-06, -6.4564716e-08, 0.00086851855, -2.4361538e-05, -3.574701e-06, -6.868703e-08, 0.0008801366, -2.2111624e-05, -3.5515584e-06, -7.2679036e-08, 0.0008906312, -1.9868156e-05, -3.5252497e-06, -7.6539024e-08, 0.0009000062, -1.76333e-05, -3.4958457e-06, -8.026543e-08, 0.00090826635, -1.5409183e-05, -3.4634188e-06, -8.385681e-08, 0.0009154175, -1.3197895e-05, -3.4280433e-06, -8.7311875e-08, 0.00092146674, -1.1001483e-05, -3.3897954e-06, -9.0629456e-08, 0.00092642184, -8.82195e-06, -3.3487527e-06, -9.380853e-08, 0.0009302918, -6.66126e-06, -3.3049944e-06, -9.684821e-08, 0.00093308656, -4.521327e-06, -3.258601e-06, -9.9747744e-08, 0.0009348169, -2.4040214e-06, -3.2096552e-06, -1.0250651e-07, 0.00093549467, -3.1116593e-07, -3.1582395e-06, -1.05124016e-07, 0.00093513244, 1.7554657e-06, -3.104439e-06, -1.075999e-07, 0.00093374384, 3.794149e-06, -3.0483386e-06, -1.0993395e-07, 0.00093134324, 5.8032097e-06, -2.9900255e-06, -1.1212607e-07, 0.00092794583, 7.7810255e-06, -2.9295866e-06, -1.14176274e-07, 0.0009235677, 9.726027e-06, -2.8671104e-06, -1.16084735e-07, 0.0009182255, 1.16366955e-05, -2.802686e-06, -1.1785174e-07, 0.0009119369, 1.3511569e-05, -2.7364024e-06, -1.1947768e-07, 0.00090472016, 1.5349236e-05, -2.6683504e-06, -1.209631e-07, 0.00089659414, 1.7148348e-05, -2.5986199e-06, -1.2230863e-07, 0.00088757847, 1.8907602e-05, -2.527302e-06, -1.2351505e-07, 0.00087769335, 2.0625757e-05, -2.4544881e-06, -1.2458324e-07, 0.00086695974, 2.230163e-05, -2.3802693e-06, -1.2551418e-07, 0.000855399, 2.3934092e-05, -2.3047369e-06, -1.2630899e-07, 0.0008430331, 2.552207e-05, -2.2279826e-06, -1.2696887e-07, 0.0008298845, 2.7064552e-05, -2.1500975e-06, -1.2749514e-07, 0.00081597624, 2.8560584e-05, -2.071173e-06, -1.2788924e-07, 0.00080133183, 3.0009267e-05, -1.9913e-06, -1.2815268e-07, 0.000785975, 3.1409763e-05, -1.910569e-06, -1.282871e-07, 0.0007699302, 3.2761287e-05, -1.8290699e-06, -1.2829419e-07, 0.00075322203, 3.406312e-05, -1.746893e-06, -1.281758e-07, 0.00073587545, 3.531459e-05, -1.6641271e-06, -1.2793382e-07, 0.00071791594, 3.6515103e-05, -1.5808608e-06, -1.2757022e-07, 0.00069936895, 3.7664096e-05, -1.497182e-06, -1.270871e-07, 0.0006802605, 3.876108e-05, -1.4131775e-06, -1.2648664e-07, 0.0006606166, 3.9805625e-05, -1.3289335e-06, -1.2577102e-07, 0.00064046367, 4.079735e-05, -1.2445354e-06, -1.2494262e-07, 0.0006198281, 4.1735933e-05, -1.1600672e-06, -1.2400376e-07, 0.00059873663, 4.2621108e-05, -1.0756123e-06, -1.2295696e-07, 0.000577216, 4.3452666e-05, -9.912526e-07, -1.218047e-07, 0.00055529294, 4.4230455e-05, -9.070691e-07, -1.2054959e-07, 0.00053299445, 4.495437e-05, -8.231413e-07, -1.1919426e-07, 0.00051034754, 4.562437e-05, -7.3954754e-07, -1.1774143e-07, 0.0004873791, 4.6240453e-05, -6.563648e-07, -1.1619386e-07, 0.00046411608, 4.680269e-05, -5.7366873e-07, -1.14554354e-07, 0.00044058537, 4.7311183e-05, -4.915332e-07, -1.12825774e-07, 0.00041681383, 4.77661e-05, -4.100309e-07, -1.11011026e-07, 0.00039282817, 4.816765e-05, -3.292328e-07, -1.09113046e-07, 0.00036865502, 4.85161e-05, -2.4920823e-07, -1.07134824e-07, 0.00034432087, 4.8811755e-05, -1.7002498e-07, -1.0507937e-07, 0.000319852, 4.9054976e-05, -9.1749e-08, -1.0294975e-07, 0.00029527457, 4.924617e-05, -1.4444599e-08, -1.0074902e-07, 0.00027061443, 4.938578e-05, 6.182573e-08, -9.848029e-08, 0.0002458973, 4.9474307e-05, 1.3700131e-07, -9.61467e-08, 0.00022114856, 4.9512284e-05, 2.1102329e-07, -9.3751375e-08, 0.00019639333, 4.95003e-05, 2.8383474e-07, -9.129749e-08, 0.00017165647, 4.943897e-05, 3.5538062e-07, -8.8788205e-08, 0.00014696248, 4.9328963e-05, 4.256078e-07, -8.6226706e-08, 0.0001223355, 4.9170976e-05, 4.9446516e-07, -8.3616186e-08, 9.779938e-05, 4.8965747e-05, 5.619035e-07, -8.0959836e-08, 7.337751e-05, 4.8714057e-05, 6.278757e-07, -7.8260854e-08, 4.909293e-05, 4.8416714e-05, 6.923366e-07, -7.552242e-08, 2.496826e-05, 4.807457e-05, 7.5524315e-07, -7.2747724e-08, 1.0256822e-06, 4.7688496e-05, 8.1655435e-07, -6.9939944e-08, -2.2713066e-05, 4.7259407e-05, 8.762311e-07, -6.710225e-08, -4.6226713e-05, 4.6788246e-05, 9.342367e-07, -6.423778e-08, -6.949446e-05, 4.627598e-05, 9.905363e-07, -6.134968e-08, -9.249601e-05, 4.5723613e-05, 1.0450971e-06, -5.844107e-08, -0.00011521156, 4.5132165e-05, 1.0978886e-06, -5.5515038e-08, -0.00013762184, 4.4502685e-05, 1.1488822e-06, -5.2574652e-08, -0.00015970808, 4.383625e-05, 1.1980516e-06, -4.9622958e-08, -0.00018145211, 4.3133958e-05, 1.2453723e-06, -4.666296e-08, -0.00020283625, 4.239692e-05, 1.2908224e-06, -4.3697653e-08, -0.00022384342, 4.1626285e-05, 1.3343815e-06, -4.0729972e-08, -0.00024445713, 4.08232e-05, 1.3760317e-06, -3.7762828e-08, -0.00026466142, 3.998884e-05, 1.415757e-06, -3.479909e-08, -0.00028444096, 3.9124403e-05, 1.4535434e-06, -3.184159e-08, -0.000303781, 3.823108e-05, 1.4893791e-06, -2.8893115e-08, -0.00032266742, 3.7310096e-05, 1.5232544e-06, -2.5956403e-08, -0.0003410867, 3.636268e-05, 1.5551611e-06, -2.3034145e-08};
endpackage
`endif
