`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam N = 4;
	localparam M = 4;
	localparam real Lfr[0:3] = {0.99237525, 0.99237525, 0.98275226, 0.98275226};
	localparam real Lfi[0:3] = {0.034385014, -0.034385014, 0.013845935, -0.013845935};
	localparam real Lbr[0:3] = {0.99237525, 0.99237525, 0.98275226, 0.98275226};
	localparam real Lbi[0:3] = {0.034385014, -0.034385014, 0.013845935, -0.013845935};
	localparam real Wfr[0:3] = {-3.445485e-06, -3.445485e-06, 1.0250402e-06, 1.0250402e-06};
	localparam real Wfi[0:3] = {-1.3232673e-07, 1.3232673e-07, 1.9739732e-06, -1.9739732e-06};
	localparam real Wbr[0:3] = {3.445485e-06, 3.445485e-06, -1.0250402e-06, -1.0250402e-06};
	localparam real Wbi[0:3] = {1.3232673e-07, -1.3232673e-07, -1.9739732e-06, 1.9739732e-06};
	localparam real Ffr[0:3][0:99] = '{
		'{-499.3932, -35.12005, 2.7881117, -0.020694872, -516.5158, -33.36749, 2.800282, -0.025561018, -532.7579, -31.598091, 2.808808, -0.030327287, -548.1115, -29.814283, 2.8137302, -0.034989163, -562.5702, -28.018482, 2.8150935, -0.039542332, -576.1284, -26.213083, 2.8129454, -0.043982662, -588.78204, -24.40046, 2.807338, -0.04830623, -600.5281, -22.58296, 2.798327, -0.052509304, -611.36456, -20.762909, 2.7859707, -0.056588367, -621.2909, -18.942598, 2.7703316, -0.060540088, -630.3075, -17.12429, 2.7514753, -0.06436135, -638.4159, -15.310215, 2.72947, -0.068049245, -645.6188, -13.502561, 2.7043872, -0.071601056, -651.9199, -11.703479, 2.676301, -0.0750143, -657.32404, -9.915084, 2.6452882, -0.07828667, -661.8371, -8.139442, 2.6114287, -0.081416085, -665.46594, -6.3785796, 2.5748043, -0.08440067, -668.21844, -4.6344724, 2.5354989, -0.08723875, -670.1035, -2.9090493, 2.4935987, -0.08992885, -671.1309, -1.2041888, 2.4491925, -0.092469715, -671.31146, 0.4782819, 2.4023702, -0.09486028, -670.6567, 2.1365898, 2.3532236, -0.09709968, -669.1792, 3.7690158, 2.3018465, -0.099187255, -666.8923, 5.373898, 2.248334, -0.10112256, -663.8101, 6.9496317, 2.192782, -0.1029053},
		'{-499.3932, -35.12005, 2.7881117, -0.020694872, -516.5158, -33.36749, 2.800282, -0.025561018, -532.7579, -31.598091, 2.808808, -0.030327287, -548.1115, -29.814283, 2.8137302, -0.034989163, -562.5702, -28.018482, 2.8150935, -0.039542332, -576.1284, -26.213083, 2.8129454, -0.043982662, -588.78204, -24.40046, 2.807338, -0.04830623, -600.5281, -22.58296, 2.798327, -0.052509304, -611.36456, -20.762909, 2.7859707, -0.056588367, -621.2909, -18.942598, 2.7703316, -0.060540088, -630.3075, -17.12429, 2.7514753, -0.06436135, -638.4159, -15.310215, 2.72947, -0.068049245, -645.6188, -13.502561, 2.7043872, -0.071601056, -651.9199, -11.703479, 2.676301, -0.0750143, -657.32404, -9.915084, 2.6452882, -0.07828667, -661.8371, -8.139442, 2.6114287, -0.081416085, -665.46594, -6.3785796, 2.5748043, -0.08440067, -668.21844, -4.6344724, 2.5354989, -0.08723875, -670.1035, -2.9090493, 2.4935987, -0.08992885, -671.1309, -1.2041888, 2.4491925, -0.092469715, -671.31146, 0.4782819, 2.4023702, -0.09486028, -670.6567, 2.1365898, 2.3532236, -0.09709968, -669.1792, 3.7690158, 2.3018465, -0.099187255, -666.8923, 5.373898, 2.248334, -0.10112256, -663.8101, 6.9496317, 2.192782, -0.1029053},
		'{497.6496, 35.007595, -2.7170272, 0.2651753, 514.7302, 33.321728, -2.6104865, 0.25808808, 530.97815, 31.676888, -2.506292, 0.2511156, 546.4138, 30.072489, -2.404415, 0.24425738, 561.0573, 28.507938, -2.3048258, 0.23751289, 574.9283, 26.982645, -2.207496, 0.23088157, 588.0464, 25.496023, -2.112396, 0.2243628, 600.43066, 24.047482, -2.0194967, 0.21795596, 612.1001, 22.636436, -1.9287685, 0.21166039, 623.07324, 21.262302, -1.8401822, 0.20547533, 633.36847, 19.924496, -1.7537081, 0.19940011, 643.0037, 18.622437, -1.6693169, 0.19343393, 651.99677, 17.355545, -1.5869788, 0.18757601, 660.365, 16.123247, -1.5066644, 0.18182553, 668.1257, 14.924966, -1.4283441, 0.17618166, 675.29553, 13.760133, -1.3519886, 0.17064354, 681.8913, 12.6281805, -1.2775682, 0.16521026, 687.92914, 11.528543, -1.2050536, 0.15988094, 693.4251, 10.460662, -1.1344154, 0.15465462, 698.39496, 9.423978, -1.0656244, 0.14953038, 702.8542, 8.417937, -0.99865144, 0.14450724, 706.81793, 7.4419904, -0.93346745, 0.13958423, 710.3011, 6.495591, -0.87004346, 0.13476035, 713.31836, 5.578198, -0.8083507, 0.1300346, 715.88403, 4.689273, -0.74836046, 0.12540592},
		'{497.6496, 35.007595, -2.7170272, 0.2651753, 514.7302, 33.321728, -2.6104865, 0.25808808, 530.97815, 31.676888, -2.506292, 0.2511156, 546.4138, 30.072489, -2.404415, 0.24425738, 561.0573, 28.507938, -2.3048258, 0.23751289, 574.9283, 26.982645, -2.207496, 0.23088157, 588.0464, 25.496023, -2.112396, 0.2243628, 600.43066, 24.047482, -2.0194967, 0.21795596, 612.1001, 22.636436, -1.9287685, 0.21166039, 623.07324, 21.262302, -1.8401822, 0.20547533, 633.36847, 19.924496, -1.7537081, 0.19940011, 643.0037, 18.622437, -1.6693169, 0.19343393, 651.99677, 17.355545, -1.5869788, 0.18757601, 660.365, 16.123247, -1.5066644, 0.18182553, 668.1257, 14.924966, -1.4283441, 0.17618166, 675.29553, 13.760133, -1.3519886, 0.17064354, 681.8913, 12.6281805, -1.2775682, 0.16521026, 687.92914, 11.528543, -1.2050536, 0.15988094, 693.4251, 10.460662, -1.1344154, 0.15465462, 698.39496, 9.423978, -1.0656244, 0.14953038, 702.8542, 8.417937, -0.99865144, 0.14450724, 706.81793, 7.4419904, -0.93346745, 0.13958423, 710.3011, 6.495591, -0.87004346, 0.13476035, 713.31836, 5.578198, -0.8083507, 0.1300346, 715.88403, 4.689273, -0.74836046, 0.12540592}};
	localparam real Ffi[0:3][0:99] = '{
		'{608.7061, -43.180954, -0.9721893, 0.14610837, 586.8933, -44.059315, -0.8689074, 0.14428274, 564.65796, -44.870716, -0.7659945, 0.1423037, 542.03375, -45.615093, -0.6635731, 0.14017588, 519.0541, -46.292454, -0.56176335, 0.13790397, 495.75244, -46.902905, -0.46068305, 0.13549283, 472.1623, -47.446617, -0.36044732, 0.1329474, 448.3169, -47.923862, -0.26116866, 0.1302727, 424.24945, -48.334972, -0.1629568, 0.12747388, 399.9929, -48.680363, -0.06591867, 0.12455613, 375.57996, -48.96053, 0.029841831, 0.12152475, 351.04312, -49.17604, 0.12422381, 0.11838509, 326.41458, -49.327526, 0.2171295, 0.11514257, 301.72617, -49.415703, 0.30846432, 0.11180263, 277.0093, -49.44135, 0.39813703, 0.1083708, 252.29509, -49.4053, 0.4860596, 0.10485262, 227.61414, -49.308475, 0.57214755, 0.10125365, 202.99658, -49.15184, 0.65631974, 0.0975795, 178.47209, -48.936428, 0.7384987, 0.09383578, 154.06978, -48.663326, 0.81861025, 0.09002811, 129.81819, -48.33369, 0.8965841, 0.08616209, 105.74531, -47.94871, 0.9723534, 0.08224336, 81.878494, -47.50965, 1.0458552, 0.078277506, 58.244457, -47.017807, 1.1170298, 0.07427011, 34.869263, -46.474525, 1.1858218, 0.070226714},
		'{-608.7061, 43.180954, 0.9721893, -0.14610837, -586.8933, 44.059315, 0.8689074, -0.14428274, -564.65796, 44.870716, 0.7659945, -0.1423037, -542.03375, 45.615093, 0.6635731, -0.14017588, -519.0541, 46.292454, 0.56176335, -0.13790397, -495.75244, 46.902905, 0.46068305, -0.13549283, -472.1623, 47.446617, 0.36044732, -0.1329474, -448.3169, 47.923862, 0.26116866, -0.1302727, -424.24945, 48.334972, 0.1629568, -0.12747388, -399.9929, 48.680363, 0.06591867, -0.12455613, -375.57996, 48.96053, -0.029841831, -0.12152475, -351.04312, 49.17604, -0.12422381, -0.11838509, -326.41458, 49.327526, -0.2171295, -0.11514257, -301.72617, 49.415703, -0.30846432, -0.11180263, -277.0093, 49.44135, -0.39813703, -0.1083708, -252.29509, 49.4053, -0.4860596, -0.10485262, -227.61414, 49.308475, -0.57214755, -0.10125365, -202.99658, 49.15184, -0.65631974, -0.0975795, -178.47209, 48.936428, -0.7384987, -0.09383578, -154.06978, 48.663326, -0.81861025, -0.09002811, -129.81819, 48.33369, -0.8965841, -0.08616209, -105.74531, 47.94871, -0.9723534, -0.08224336, -81.878494, 47.50965, -1.0458552, -0.078277506, -58.244457, 47.017807, -1.1170298, -0.07427011, -34.869263, 46.474525, -1.1858218, -0.070226714},
		'{-1853.5363, 78.15038, -4.3101377, 0.18153787, -1814.6765, 77.28718, -4.2734175, 0.18207835, -1776.2505, 76.41552, -4.235855, 0.18251137, -1738.2623, 75.53612, -4.197498, 0.18284039, -1700.7156, 74.64967, -4.158392, 0.18306878, -1663.6136, 73.75685, -4.118582, 0.18319984, -1626.9597, 72.858315, -4.07811, 0.18323682, -1590.7562, 71.95469, -4.03702, 0.18318291, -1555.0057, 71.04659, -3.9953523, 0.18304123, -1519.7102, 70.13462, -3.9531472, 0.1828148, -1484.8717, 69.21935, -3.9104433, 0.18250667, -1450.4913, 68.301346, -3.8672786, 0.18211971, -1416.5707, 67.38115, -3.82369, 0.18165684, -1383.1105, 66.459274, -3.7797132, 0.18112083, -1350.1116, 65.53625, -3.7353828, 0.18051444, -1317.5743, 64.61254, -3.6907325, 0.17984039, -1285.499, 63.688644, -3.6457953, 0.17910126, -1253.8856, 62.765007, -3.6006026, 0.17829965, -1222.7339, 61.842075, -3.5551853, 0.17743808, -1192.0435, 60.920277, -3.5095735, 0.17651902, -1161.8134, 60.000023, -3.4637957, 0.17554484, -1132.0431, 59.08171, -3.4178803, 0.17451793, -1102.7313, 58.165726, -3.3718543, 0.17344056, -1073.8768, 57.252434, -3.325744, 0.17231499, -1045.4784, 56.342194, -3.2795746, 0.1711434},
		'{1853.5363, -78.15038, 4.3101377, -0.18153787, 1814.6765, -77.28718, 4.2734175, -0.18207835, 1776.2505, -76.41552, 4.235855, -0.18251137, 1738.2623, -75.53612, 4.197498, -0.18284039, 1700.7156, -74.64967, 4.158392, -0.18306878, 1663.6136, -73.75685, 4.118582, -0.18319984, 1626.9597, -72.858315, 4.07811, -0.18323682, 1590.7562, -71.95469, 4.03702, -0.18318291, 1555.0057, -71.04659, 3.9953523, -0.18304123, 1519.7102, -70.13462, 3.9531472, -0.1828148, 1484.8717, -69.21935, 3.9104433, -0.18250667, 1450.4913, -68.301346, 3.8672786, -0.18211971, 1416.5707, -67.38115, 3.82369, -0.18165684, 1383.1105, -66.459274, 3.7797132, -0.18112083, 1350.1116, -65.53625, 3.7353828, -0.18051444, 1317.5743, -64.61254, 3.6907325, -0.17984039, 1285.499, -63.688644, 3.6457953, -0.17910126, 1253.8856, -62.765007, 3.6006026, -0.17829965, 1222.7339, -61.842075, 3.5551853, -0.17743808, 1192.0435, -60.920277, 3.5095735, -0.17651902, 1161.8134, -60.000023, 3.4637957, -0.17554484, 1132.0431, -59.08171, 3.4178803, -0.17451793, 1102.7313, -58.165726, 3.3718543, -0.17344056, 1073.8768, -57.252434, 3.325744, -0.17231499, 1045.4784, -56.342194, 3.2795746, -0.1711434}};
	localparam real Fbr[0:3][0:99] = '{
		'{499.3932, -35.12005, -2.7881117, -0.020694872, 516.5158, -33.36749, -2.800282, -0.025561018, 532.7579, -31.598091, -2.808808, -0.030327287, 548.1115, -29.814283, -2.8137302, -0.034989163, 562.5702, -28.018482, -2.8150935, -0.039542332, 576.1284, -26.213083, -2.8129454, -0.043982662, 588.78204, -24.40046, -2.807338, -0.04830623, 600.5281, -22.58296, -2.798327, -0.052509304, 611.36456, -20.762909, -2.7859707, -0.056588367, 621.2909, -18.942598, -2.7703316, -0.060540088, 630.3075, -17.12429, -2.7514753, -0.06436135, 638.4159, -15.310215, -2.72947, -0.068049245, 645.6188, -13.502561, -2.7043872, -0.071601056, 651.9199, -11.703479, -2.676301, -0.0750143, 657.32404, -9.915084, -2.6452882, -0.07828667, 661.8371, -8.139442, -2.6114287, -0.081416085, 665.46594, -6.3785796, -2.5748043, -0.08440067, 668.21844, -4.6344724, -2.5354989, -0.08723875, 670.1035, -2.9090493, -2.4935987, -0.08992885, 671.1309, -1.2041888, -2.4491925, -0.092469715, 671.31146, 0.4782819, -2.4023702, -0.09486028, 670.6567, 2.1365898, -2.3532236, -0.09709968, 669.1792, 3.7690158, -2.3018465, -0.099187255, 666.8923, 5.373898, -2.248334, -0.10112256, 663.8101, 6.9496317, -2.192782, -0.1029053},
		'{499.3932, -35.12005, -2.7881117, -0.020694872, 516.5158, -33.36749, -2.800282, -0.025561018, 532.7579, -31.598091, -2.808808, -0.030327287, 548.1115, -29.814283, -2.8137302, -0.034989163, 562.5702, -28.018482, -2.8150935, -0.039542332, 576.1284, -26.213083, -2.8129454, -0.043982662, 588.78204, -24.40046, -2.807338, -0.04830623, 600.5281, -22.58296, -2.798327, -0.052509304, 611.36456, -20.762909, -2.7859707, -0.056588367, 621.2909, -18.942598, -2.7703316, -0.060540088, 630.3075, -17.12429, -2.7514753, -0.06436135, 638.4159, -15.310215, -2.72947, -0.068049245, 645.6188, -13.502561, -2.7043872, -0.071601056, 651.9199, -11.703479, -2.676301, -0.0750143, 657.32404, -9.915084, -2.6452882, -0.07828667, 661.8371, -8.139442, -2.6114287, -0.081416085, 665.46594, -6.3785796, -2.5748043, -0.08440067, 668.21844, -4.6344724, -2.5354989, -0.08723875, 670.1035, -2.9090493, -2.4935987, -0.08992885, 671.1309, -1.2041888, -2.4491925, -0.092469715, 671.31146, 0.4782819, -2.4023702, -0.09486028, 670.6567, 2.1365898, -2.3532236, -0.09709968, 669.1792, 3.7690158, -2.3018465, -0.099187255, 666.8923, 5.373898, -2.248334, -0.10112256, 663.8101, 6.9496317, -2.192782, -0.1029053},
		'{-497.6496, 35.007595, 2.7170272, 0.2651753, -514.7302, 33.321728, 2.6104865, 0.25808808, -530.97815, 31.676888, 2.506292, 0.2511156, -546.4138, 30.072489, 2.404415, 0.24425738, -561.0573, 28.507938, 2.3048258, 0.23751289, -574.9283, 26.982645, 2.207496, 0.23088157, -588.0464, 25.496023, 2.112396, 0.2243628, -600.43066, 24.047482, 2.0194967, 0.21795596, -612.1001, 22.636436, 1.9287685, 0.21166039, -623.07324, 21.262302, 1.8401822, 0.20547533, -633.36847, 19.924496, 1.7537081, 0.19940011, -643.0037, 18.622437, 1.6693169, 0.19343393, -651.99677, 17.355545, 1.5869788, 0.18757601, -660.365, 16.123247, 1.5066644, 0.18182553, -668.1257, 14.924966, 1.4283441, 0.17618166, -675.29553, 13.760133, 1.3519886, 0.17064354, -681.8913, 12.6281805, 1.2775682, 0.16521026, -687.92914, 11.528543, 1.2050536, 0.15988094, -693.4251, 10.460662, 1.1344154, 0.15465462, -698.39496, 9.423978, 1.0656244, 0.14953038, -702.8542, 8.417937, 0.99865144, 0.14450724, -706.81793, 7.4419904, 0.93346745, 0.13958423, -710.3011, 6.495591, 0.87004346, 0.13476035, -713.31836, 5.578198, 0.8083507, 0.1300346, -715.88403, 4.689273, 0.74836046, 0.12540592},
		'{-497.6496, 35.007595, 2.7170272, 0.2651753, -514.7302, 33.321728, 2.6104865, 0.25808808, -530.97815, 31.676888, 2.506292, 0.2511156, -546.4138, 30.072489, 2.404415, 0.24425738, -561.0573, 28.507938, 2.3048258, 0.23751289, -574.9283, 26.982645, 2.207496, 0.23088157, -588.0464, 25.496023, 2.112396, 0.2243628, -600.43066, 24.047482, 2.0194967, 0.21795596, -612.1001, 22.636436, 1.9287685, 0.21166039, -623.07324, 21.262302, 1.8401822, 0.20547533, -633.36847, 19.924496, 1.7537081, 0.19940011, -643.0037, 18.622437, 1.6693169, 0.19343393, -651.99677, 17.355545, 1.5869788, 0.18757601, -660.365, 16.123247, 1.5066644, 0.18182553, -668.1257, 14.924966, 1.4283441, 0.17618166, -675.29553, 13.760133, 1.3519886, 0.17064354, -681.8913, 12.6281805, 1.2775682, 0.16521026, -687.92914, 11.528543, 1.2050536, 0.15988094, -693.4251, 10.460662, 1.1344154, 0.15465462, -698.39496, 9.423978, 1.0656244, 0.14953038, -702.8542, 8.417937, 0.99865144, 0.14450724, -706.81793, 7.4419904, 0.93346745, 0.13958423, -710.3011, 6.495591, 0.87004346, 0.13476035, -713.31836, 5.578198, 0.8083507, 0.1300346, -715.88403, 4.689273, 0.74836046, 0.12540592}};
	localparam real Fbi[0:3][0:99] = '{
		'{-608.7061, -43.180954, 0.9721893, 0.14610837, -586.8933, -44.059315, 0.8689074, 0.14428274, -564.65796, -44.870716, 0.7659945, 0.1423037, -542.03375, -45.615093, 0.6635731, 0.14017588, -519.0541, -46.292454, 0.56176335, 0.13790397, -495.75244, -46.902905, 0.46068305, 0.13549283, -472.1623, -47.446617, 0.36044732, 0.1329474, -448.3169, -47.923862, 0.26116866, 0.1302727, -424.24945, -48.334972, 0.1629568, 0.12747388, -399.9929, -48.680363, 0.06591867, 0.12455613, -375.57996, -48.96053, -0.029841831, 0.12152475, -351.04312, -49.17604, -0.12422381, 0.11838509, -326.41458, -49.327526, -0.2171295, 0.11514257, -301.72617, -49.415703, -0.30846432, 0.11180263, -277.0093, -49.44135, -0.39813703, 0.1083708, -252.29509, -49.4053, -0.4860596, 0.10485262, -227.61414, -49.308475, -0.57214755, 0.10125365, -202.99658, -49.15184, -0.65631974, 0.0975795, -178.47209, -48.936428, -0.7384987, 0.09383578, -154.06978, -48.663326, -0.81861025, 0.09002811, -129.81819, -48.33369, -0.8965841, 0.08616209, -105.74531, -47.94871, -0.9723534, 0.08224336, -81.878494, -47.50965, -1.0458552, 0.078277506, -58.244457, -47.017807, -1.1170298, 0.07427011, -34.869263, -46.474525, -1.1858218, 0.070226714},
		'{608.7061, 43.180954, -0.9721893, -0.14610837, 586.8933, 44.059315, -0.8689074, -0.14428274, 564.65796, 44.870716, -0.7659945, -0.1423037, 542.03375, 45.615093, -0.6635731, -0.14017588, 519.0541, 46.292454, -0.56176335, -0.13790397, 495.75244, 46.902905, -0.46068305, -0.13549283, 472.1623, 47.446617, -0.36044732, -0.1329474, 448.3169, 47.923862, -0.26116866, -0.1302727, 424.24945, 48.334972, -0.1629568, -0.12747388, 399.9929, 48.680363, -0.06591867, -0.12455613, 375.57996, 48.96053, 0.029841831, -0.12152475, 351.04312, 49.17604, 0.12422381, -0.11838509, 326.41458, 49.327526, 0.2171295, -0.11514257, 301.72617, 49.415703, 0.30846432, -0.11180263, 277.0093, 49.44135, 0.39813703, -0.1083708, 252.29509, 49.4053, 0.4860596, -0.10485262, 227.61414, 49.308475, 0.57214755, -0.10125365, 202.99658, 49.15184, 0.65631974, -0.0975795, 178.47209, 48.936428, 0.7384987, -0.09383578, 154.06978, 48.663326, 0.81861025, -0.09002811, 129.81819, 48.33369, 0.8965841, -0.08616209, 105.74531, 47.94871, 0.9723534, -0.08224336, 81.878494, 47.50965, 1.0458552, -0.078277506, 58.244457, 47.017807, 1.1170298, -0.07427011, 34.869263, 46.474525, 1.1858218, -0.070226714},
		'{1853.5363, 78.15038, 4.3101377, 0.18153787, 1814.6765, 77.28718, 4.2734175, 0.18207835, 1776.2505, 76.41552, 4.235855, 0.18251137, 1738.2623, 75.53612, 4.197498, 0.18284039, 1700.7156, 74.64967, 4.158392, 0.18306878, 1663.6136, 73.75685, 4.118582, 0.18319984, 1626.9597, 72.858315, 4.07811, 0.18323682, 1590.7562, 71.95469, 4.03702, 0.18318291, 1555.0057, 71.04659, 3.9953523, 0.18304123, 1519.7102, 70.13462, 3.9531472, 0.1828148, 1484.8717, 69.21935, 3.9104433, 0.18250667, 1450.4913, 68.301346, 3.8672786, 0.18211971, 1416.5707, 67.38115, 3.82369, 0.18165684, 1383.1105, 66.459274, 3.7797132, 0.18112083, 1350.1116, 65.53625, 3.7353828, 0.18051444, 1317.5743, 64.61254, 3.6907325, 0.17984039, 1285.499, 63.688644, 3.6457953, 0.17910126, 1253.8856, 62.765007, 3.6006026, 0.17829965, 1222.7339, 61.842075, 3.5551853, 0.17743808, 1192.0435, 60.920277, 3.5095735, 0.17651902, 1161.8134, 60.000023, 3.4637957, 0.17554484, 1132.0431, 59.08171, 3.4178803, 0.17451793, 1102.7313, 58.165726, 3.3718543, 0.17344056, 1073.8768, 57.252434, 3.325744, 0.17231499, 1045.4784, 56.342194, 3.2795746, 0.1711434},
		'{-1853.5363, -78.15038, -4.3101377, -0.18153787, -1814.6765, -77.28718, -4.2734175, -0.18207835, -1776.2505, -76.41552, -4.235855, -0.18251137, -1738.2623, -75.53612, -4.197498, -0.18284039, -1700.7156, -74.64967, -4.158392, -0.18306878, -1663.6136, -73.75685, -4.118582, -0.18319984, -1626.9597, -72.858315, -4.07811, -0.18323682, -1590.7562, -71.95469, -4.03702, -0.18318291, -1555.0057, -71.04659, -3.9953523, -0.18304123, -1519.7102, -70.13462, -3.9531472, -0.1828148, -1484.8717, -69.21935, -3.9104433, -0.18250667, -1450.4913, -68.301346, -3.8672786, -0.18211971, -1416.5707, -67.38115, -3.82369, -0.18165684, -1383.1105, -66.459274, -3.7797132, -0.18112083, -1350.1116, -65.53625, -3.7353828, -0.18051444, -1317.5743, -64.61254, -3.6907325, -0.17984039, -1285.499, -63.688644, -3.6457953, -0.17910126, -1253.8856, -62.765007, -3.6006026, -0.17829965, -1222.7339, -61.842075, -3.5551853, -0.17743808, -1192.0435, -60.920277, -3.5095735, -0.17651902, -1161.8134, -60.000023, -3.4637957, -0.17554484, -1132.0431, -59.08171, -3.4178803, -0.17451793, -1102.7313, -58.165726, -3.3718543, -0.17344056, -1073.8768, -57.252434, -3.325744, -0.17231499, -1045.4784, -56.342194, -3.2795746, -0.1711434}};
	localparam real hf[0:1199] = {0.011940284, -6.1819783e-06, -8.024018e-06, 8.204753e-09, 0.0119341025, -1.8539538e-05, -8.007101e-06, 2.4590857e-08, 0.011921748, -3.087793e-05, -7.9733045e-06, 4.0907583e-08, 0.01190323, -4.3184416e-05, -7.922693e-06, 5.711045e-08, 0.011878571, -5.5446304e-05, -7.855365e-06, 7.315652e-08, 0.011847793, -6.765098e-05, -7.771447e-06, 8.9004416e-08, 0.01181093, -7.9785925e-05, -7.671095e-06, 1.0461433e-07, 0.011768021, -9.183872e-05, -7.554496e-06, 1.1994803e-07, 0.011719108, -0.00010379708, -7.4218597e-06, 1.349689e-07, 0.011664242, -0.00011564886, -7.273425e-06, 1.4964193e-07, 0.011603478, -0.00012738208, -7.109457e-06, 1.6393372e-07, 0.011536881, -0.00013898496, -6.930243e-06, 1.7781245e-07, 0.011464518, -0.00015044588, -6.7360957e-06, 1.91248e-07, 0.011386461, -0.00016175344, -6.52735e-06, 2.042118e-07, 0.011302792, -0.0001728965, -6.304362e-06, 2.1667695e-07, 0.011213593, -0.00018386412, -6.0675097e-06, 2.2861816e-07, 0.011118958, -0.00019464563, -5.8171895e-06, 2.4001173e-07, 0.01101898, -0.00020523065, -5.5538176e-06, 2.5083557e-07, 0.010913762, -0.00021560903, -5.2778278e-06, 2.6106926e-07, 0.010803408, -0.00022577097, -4.98967e-06, 2.7069387e-07, 0.010688028, -0.00023570693, -4.6898103e-06, 2.7969216e-07, 0.01056774, -0.00024540772, -4.3787304e-06, 2.8804834e-07, 0.010442661, -0.00025486446, -4.0569244e-06, 2.9574826e-07, 0.010312918, -0.0002640686, -3.7248994e-06, 3.027793e-07, 0.010178637, -0.00027301194, -3.383175e-06, 3.0913034e-07, 0.010039951, -0.00028168663, -3.032281e-06, 3.1479172e-07, 0.0098969955, -0.00029008518, -2.672757e-06, 3.1975532e-07, 0.009749913, -0.00029820052, -2.3051512e-06, 3.2401448e-07, 0.009598844, -0.00030602588, -1.93002e-06, 3.2756392e-07, 0.009443936, -0.0003135549, -1.5479261e-06, 3.303998e-07, 0.009285339, -0.00032078158, -1.1594383e-06, 3.325197e-07, 0.009123205, -0.0003277004, -7.6513027e-07, 3.3392251e-07, 0.008957691, -0.00033430613, -3.6557958e-07, 3.3460844e-07, 0.008788953, -0.000340594, 3.863335e-08, 3.3457906e-07, 0.008617151, -0.00034655962, 4.469259e-07, 3.338371e-07, 0.0084424475, -0.00035219904, 8.587143e-07, 3.323867e-07, 0.008265006, -0.00035750863, 1.2734147e-06, 3.3023298e-07, 0.008084994, -0.00036248527, 1.6904436e-06, 3.2738242e-07, 0.0079025775, -0.0003671262, 2.1092192e-06, 3.2384258e-07, 0.007717924, -0.00037142902, 2.529162e-06, 3.1962207e-07, 0.0075312047, -0.00037539183, 2.9496955e-06, 3.1473067e-07, 0.007342589, -0.0003790131, 3.3702477e-06, 3.0917906e-07, 0.0071522486, -0.00038229168, 3.7902503e-06, 3.0297903e-07, 0.0069603547, -0.00038522683, 4.2091415e-06, 2.9614327e-07, 0.0067670792, -0.0003878182, 4.626366e-06, 2.886854e-07, 0.006572594, -0.00039006592, 5.0413737e-06, 2.8061996e-07, 0.0063770707, -0.0003919704, 5.4536245e-06, 2.7196222e-07, 0.006180681, -0.0003935325, 5.8625856e-06, 2.6272835e-07, 0.005983595, -0.00039475344, 6.267733e-06, 2.529353e-07, 0.0057859835, -0.00039563482, 6.668553e-06, 2.4260066e-07, 0.0055880165, -0.00039617866, 7.0645415e-06, 2.3174275e-07, 0.005389861, -0.00039638727, 7.4552063e-06, 2.2038053e-07, 0.0051916847, -0.0003962634, 7.840066e-06, 2.0853356e-07, 0.0049936525, -0.0003958101, 8.218651e-06, 1.9622199e-07, 0.004795929, -0.00039503071, 8.590505e-06, 1.8346643e-07, 0.0045986753, -0.00039392908, 8.955183e-06, 1.7028802e-07, 0.0044020526, -0.00039250925, 9.312257e-06, 1.5670835e-07, 0.0042062183, -0.00039077562, 9.6613085e-06, 1.4274937e-07, 0.004011329, -0.0003887329, 1.0001936e-05, 1.2843343e-07, 0.0038175362, -0.00038638615, 1.0333753e-05, 1.1378318e-07, 0.0036249922, -0.00038374067, 1.0656387e-05, 9.882157e-08, 0.0034338445, -0.00038080206, 1.096948e-05, 8.3571805e-08, 0.003244238, -0.0003775762, 1.1272693e-05, 6.805727e-08, 0.0030563152, -0.00037406923, 1.15656985e-05, 5.2301523e-08, 0.0028702146, -0.00037028757, 1.1848189e-05, 3.6328274e-08, 0.0026860721, -0.00036623792, 1.2119873e-05, 2.016131e-08, 0.0025040202, -0.0003619271, 1.2380473e-05, 3.8244825e-09, 0.0023241874, -0.00035736224, 1.2629732e-05, -1.265834e-08, 0.0021466992, -0.0003525507, 1.2867406e-05, -2.92633e-08, 0.0019716767, -0.00034749997, 1.3093272e-05, -4.5966587e-08, 0.0017992377, -0.00034221783, 1.33071235e-05, -6.274448e-08, 0.0016294961, -0.0003367121, 1.35087685e-05, -7.957337e-08, 0.0014625615, -0.00033099094, 1.3698036e-05, -9.6429794e-08, 0.0012985397, -0.00032506252, 1.387477e-05, -1.13290476e-07, 0.0011375322, -0.00031893523, 1.4038833e-05, -1.3013234e-07, 0.0009796362, -0.00031261757, 1.4190105e-05, -1.4693258e-07, 0.0008249449, -0.0003061182, 1.43284815e-05, -1.6366863e-07, 0.00067354686, -0.00029944582, 1.4453879e-05, -1.8031824e-07, 0.0005255264, -0.00029260933, 1.4566228e-05, -1.9685949e-07, 0.0003809634, -0.0002856176, 1.46654775e-05, -2.1327081e-07, 0.00023993319, -0.00027847965, 1.4751593e-05, -2.2953101e-07, 0.00010250661, -0.00027120457, 1.4824558e-05, -2.4561933e-07, -3.1250034e-05, -0.00026380146, 1.488437e-05, -2.615154e-07, -0.00016127502, -0.00025627948, 1.4931046e-05, -2.7719932e-07, -0.00028751124, -0.00024864782, 1.4964618e-05, -2.926517e-07, -0.0004099061, -0.00024091572, 1.4985132e-05, -3.0785355e-07, -0.0005284117, -0.00023309235, 1.49926545e-05, -3.2278655e-07, -0.00064298476, -0.00022518694, 1.4987263e-05, -3.374328e-07, -0.00075358653, -0.00021720871, 1.4969053e-05, -3.5177496e-07, -0.00086018286, -0.00020916681, 1.4938134e-05, -3.6579627e-07, -0.00096274423, -0.00020107039, 1.4894629e-05, -3.794806e-07, -0.0010612457, -0.00019292852, 1.4838679e-05, -3.9281244e-07, -0.0011556667, -0.00018475026, 1.4770433e-05, -4.0577677e-07, -0.0012459913, -0.00017654453, 1.469006e-05, -4.183593e-07, -0.0013322082, -0.00016832027, 1.4597737e-05, -4.3054638e-07, -0.00141431, -0.00016008626, 1.4493659e-05, -4.42325e-07, -0.0014922943, -0.0001518512, 1.4378028e-05, -4.5368273e-07, -0.0015661624, -0.0001436237, 1.4251062e-05, -4.6460795e-07, -0.0016359206, -0.00013541225, 1.41129885e-05, -4.7508965e-07, -0.0017015787, -0.00012722521, 1.3964048e-05, -4.851175e-07, -0.0017631513, -0.00011907082, 1.3804491e-05, -4.946818e-07, -0.0018206564, -0.00011095717, 1.3634577e-05, -5.0377366e-07, -0.0018741165, -0.00010289221, 1.3454577e-05, -5.123848e-07, -0.001923558, -9.488373e-05, 1.3264772e-05, -5.205078e-07, -0.001969011, -8.693937e-05, 1.306545e-05, -5.281357e-07, -0.0020105094, -7.906658e-05, 1.2856909e-05, -5.352623e-07, -0.0020480906, -7.1272654e-05, 1.2639454e-05, -5.4188234e-07, -0.0020817963, -6.3564694e-05, 1.2413399e-05, -5.4799096e-07, -0.0021116708, -5.594962e-05, 1.2179065e-05, -5.535842e-07, -0.0021377625, -4.8434144e-05, 1.1936777e-05, -5.5865866e-07, -0.0021601226, -4.1024792e-05, 1.1686869e-05, -5.6321176e-07, -0.002178806, -3.3727883e-05, 1.1429678e-05, -5.6724144e-07, -0.0021938703, -2.654952e-05, 1.116555e-05, -5.707466e-07, -0.0022053763, -1.94956e-05, 1.08948325e-05, -5.737265e-07, -0.0022133875, -1.257179e-05, 1.0617877e-05, -5.761812e-07, -0.0022179708, -5.7835446e-06, 1.033504e-05, -5.781115e-07, -0.0022191945, 8.6391225e-07, 1.0046682e-05, -5.795188e-07, -0.002217131, 7.365586e-06, 9.753164e-06, -5.8040507e-07, -0.002211854, 1.3716714e-05, 9.45485e-06, -5.80773e-07, -0.0022034403, 1.991277e-05, 9.152107e-06, -5.806259e-07, -0.0021919678, 2.5949465e-05, 8.845302e-06, -5.799676e-07, -0.0021775179, 3.1822747e-05, 8.534802e-06, -5.7880266e-07, -0.002160173, 3.7528807e-05, 8.220977e-06, -5.7713606e-07, -0.0021400177, 4.3064083e-05, 7.904194e-06, -5.7497346e-07, -0.002117138, 4.8425245e-05, 7.58482e-06, -5.7232114e-07, -0.002091622, 5.3609227e-05, 7.263224e-06, -5.691858e-07, -0.0020635587, 5.8613183e-05, 6.9397693e-06, -5.655747e-07, -0.0020330392, 6.3434534e-05, 6.6148195e-06, -5.614956e-07, -0.002000155, 6.8070935e-05, 6.288736e-06, -5.569569e-07, -0.0019649994, 7.2520284e-05, 5.961877e-06, -5.5196716e-07, -0.0019276662, 7.678073e-05, 5.634597e-06, -5.4653583e-07, -0.0018882505, 8.085066e-05, 5.3072476e-06, -5.406724e-07, -0.0018468476, 8.472871e-05, 4.980177e-06, -5.34387e-07, -0.0018035539, 8.841373e-05, 4.6537284e-06, -5.2769025e-07, -0.0017584661, 9.190485e-05, 4.32824e-06, -5.2059295e-07, -0.0017116815, 9.5201394e-05, 4.0040454e-06, -5.131064e-07, -0.0016632973, 9.830295e-05, 3.681473e-06, -5.0524216e-07, -0.001613411, 0.00010120933, 3.360845e-06, -4.970123e-07, -0.0015621204, 0.00010392056, 3.0424783e-06, -4.88429e-07, -0.001509523, 0.0001064369, 2.7266829e-06, -4.79505e-07, -0.001455716, 0.00010875883, 2.413762e-06, -4.7025296e-07, -0.0014007965, 0.00011088706, 2.1040125e-06, -4.6068612e-07, -0.001344861, 0.0001128225, 1.7977234e-06, -4.508178e-07, -0.0012880058, 0.00011456626, 1.4951765e-06, -4.4066155e-07, -0.0012303265, 0.00011611969, 1.1966463e-06, -4.302312e-07, -0.0011719177, 0.00011748432, 9.023985e-07, -4.1954067e-07, -0.0011128733, 0.00011866187, 6.126912e-07, -4.0860408e-07, -0.0010532866, 0.000119654265, 3.2777407e-07, -3.9743568e-07, -0.0009932496, 0.000120463614, 4.7888012e-08, -3.8604986e-07, -0.00093285315, 0.0001210922, -2.2673481e-07, -3.7446114e-07, -0.0008721871, 0.00012154251, -4.958712e-07, -3.62684e-07, -0.00081133994, 0.00012181716, -7.5930694e-07, -3.5073316e-07, -0.0007503987, 0.00012191897, -1.0168372e-06, -3.386232e-07, -0.00068944925, 0.000121850906, -1.2682666e-06, -3.2636893e-07, -0.0006285756, 0.00012161609, -1.5134091e-06, -3.1398497e-07, -0.00056786044, 0.00012121779, -1.7520883e-06, -3.0148607e-07, -0.00050738454, 0.00012065941, -1.9841377e-06, -2.8888687e-07, -0.0004472271, 0.00011994451, -2.2094002e-06, -2.7620203e-07, -0.0003874655, 0.00011907677, -2.427729e-06, -2.6344605e-07, -0.00032817517, 0.000118059994, -2.6389869e-06, -2.506335e-07, -0.0002694297, 0.0001168981, -2.8430466e-06, -2.3777866e-07, -0.00021130059, 0.00011559514, -3.039791e-06, -2.2489587e-07, -0.00015385737, 0.00011415523, -3.2291125e-06, -2.1199925e-07, -9.7167474e-05, 0.000112582624, -3.4109146e-06, -1.9910277e-07, -4.129615e-05, 0.00011088165, -3.5851092e-06, -1.8622028e-07, 1.3693514e-05, 0.000109056724, -3.7516195e-06, -1.7336544e-07, 6.7740664e-05, 0.000107112355, -3.910378e-06, -1.6055168e-07, 0.00012078672, 0.0001050531, -4.0613268e-06, -1.4779228e-07, 0.00017277538, 0.0001028836, -4.2044185e-06, -1.3510027e-07, 0.00022365272, 0.00010060855, -4.3396144e-06, -1.2248844e-07, 0.00027336713, 9.823271e-05, -4.4668873e-06, -1.09969385e-07, 0.00032186942, 9.576087e-05, -4.5862175e-06, -9.755537e-08, 0.00036911282, 9.319787e-05, -4.6975956e-06, -8.525845e-08, 0.00041505293, 9.054859e-05, -4.8010224e-06, -7.309037e-08, 0.00045964782, 8.781791e-05, -4.896506e-06, -6.106258e-08, 0.0005028581, 8.501077e-05, -4.984066e-06, -4.9186248e-08, 0.0005446467, 8.21321e-05, -5.063729e-06, -3.7472216e-08, 0.0005849791, 7.9186844e-05, -5.1355314e-06, -2.593101e-08, 0.00062382326, 7.617996e-05, -5.199517e-06, -1.45728265e-08, 0.0006611496, 7.311639e-05, -5.2557402e-06, -3.4075192e-09, 0.00069693103, 7.000107e-05, -5.3042622e-06, 7.5554e-09, 0.0007311429, 6.683892e-05, -5.3451527e-06, 1.8306773e-08, 0.0007637629, 6.363485e-05, -5.3784884e-06, 2.8837803e-08, 0.00079477153, 6.039373e-05, -5.4043558e-06, 3.914006e-08, 0.0008241513, 5.712041e-05, -5.422847e-06, 4.920548e-08, 0.0008518874, 5.3819695e-05, -5.4340626e-06, 5.902638e-08, 0.0008779672, 5.0496346e-05, -5.4381094e-06, 6.859546e-08, 0.00090238074, 4.715509e-05, -5.4351017e-06, 7.79058e-08, 0.0009251201, 4.3800588e-05, -5.4251605e-06, 8.6950884e-08, 0.00094617985, 4.0437444e-05, -5.408412e-06, 9.572456e-08, 0.0009655569, 3.7070215e-05, -5.384991e-06, 1.0422109e-07, 0.0009832501, 3.3703367e-05, -5.3550352e-06, 1.1243513e-07, 0.000999261, 3.034132e-05, -5.3186905e-06, 1.2036173e-07, 0.001013593, 2.6988402e-05, -5.276107e-06, 1.2799634e-07, 0.0010262517, 2.3648865e-05, -5.22744e-06, 1.3533482e-07, 0.0010372448, 2.032688e-05, -5.17285e-06, 1.423734e-07, 0.0010465821, 1.7026527e-05, -5.112502e-06, 1.4910871e-07, 0.0010542755, 1.3751798e-05, -5.046566e-06, 1.5553783e-07, 0.0010603388, 1.050659e-05, -4.9752152e-06, 1.6165818e-07, 0.0010647877, 7.2947e-06, -4.898627e-06, 1.6746759e-07, 0.0010676397, 4.119824e-06, -4.8169827e-06, 1.7296428e-07, 0.0010689143, 9.855555e-07, -4.730466e-06, 1.7814686e-07, 0.0010686326, -2.1046212e-06, -4.639265e-06, 1.8301432e-07, 0.0010668176, -5.147331e-06, -4.5435704e-06, 1.8756604e-07, 0.0010634938, -8.139311e-06, -4.4435737e-06, 1.9180179e-07, 0.0010586872, -1.1077412e-05, -4.3394707e-06, 1.9572165e-07, 0.0010524258, -1.3958604e-05, -4.2314587e-06, 1.9932614e-07, 0.0010447387, -1.6779974e-05, -4.119736e-06, 2.026161e-07, 0.0010356563, -1.953873e-05, -4.0045024e-06, 2.0559277e-07, 0.0010252108, -2.2232203e-05, -3.8859603e-06, 2.0825766e-07, 0.0010134354, -2.4857845e-05, -3.7643117e-06, 2.1061268e-07, 0.0010003647, -2.741324e-05, -3.6397594e-06, 2.1266008e-07, 0.0009860343, -2.989609e-05, -3.512507e-06, 2.1440243e-07, 0.000970481, -3.230423e-05, -3.3827585e-06, 2.1584259e-07, 0.0009537428, -3.4635617e-05, -3.2507169e-06, 2.1698379e-07, 0.0009358585, -3.6888345e-05, -3.116586e-06, 2.1782952e-07, 0.00091686787, -3.906063e-05, -2.9805683e-06, 2.1838359e-07, 0.00089681154, -4.1150815e-05, -2.842866e-06, 2.1865007e-07, 0.000875731, -4.3157386e-05, -2.7036797e-06, 2.1863337e-07, 0.0008536683, -4.5078945e-05, -2.5632094e-06, 2.1833812e-07, 0.00083066645, -4.691423e-05, -2.421653e-06, 2.177692e-07, 0.00080676866, -4.86621e-05, -2.2792071e-06, 2.1693181e-07, 0.00078201905, -5.0321552e-05, -2.1360665e-06, 2.1583132e-07, 0.000756462, -5.1891704e-05, -1.9924237e-06, 2.1447337e-07, 0.00073014235, -5.337181e-05, -1.8484684e-06, 2.1286382e-07, 0.0007031053, -5.4761233e-05, -1.7043886e-06, 2.1100877e-07, 0.00067539635, -5.6059478e-05, -1.5603694e-06, 2.0891444e-07, 0.0006470611, -5.7266167e-05, -1.4165925e-06, 2.0658733e-07, 0.00061814545, -5.8381043e-05, -1.273237e-06, 2.0403407e-07, 0.0005886954, -5.940397e-05, -1.1304786e-06, 2.012615e-07, 0.0005587568, -6.0334933e-05, -9.884898e-07, 1.9827658e-07, 0.0005283758, -6.117403e-05, -8.474391e-07, 1.9508646e-07, 0.0004975981, -6.192149e-05, -7.074916e-07, 1.9169838e-07, 0.0004664695, -6.257763e-05, -5.6880845e-07, 1.8811977e-07, 0.0004350356, -6.31429e-05, -4.3154677e-07, 1.8435814e-07, 0.00040334166, -6.3617845e-05, -2.958595e-07, 1.8042111e-07, 0.0003714327, -6.400313e-05, -1.6189534e-07, 1.763164e-07, 0.00033935334, -6.4299515e-05, -2.9798583e-08, 1.7205184e-07, 0.00030714786, -6.450787e-05, 1.0029098e-07, 1.6763529e-07, 0.00027485998, -6.4629145e-05, 2.2823818e-07, 1.6307472e-07, 0.00024253305, -6.466442e-05, 3.5391255e-07, 1.5837811e-07, 0.00021020972, -6.461484e-05, 4.7718845e-07, 1.5355353e-07, 0.00017793213, -6.4481654e-05, 5.979451e-07, 1.4860906e-07, 0.00014574177, -6.42662e-05, 7.1606667e-07, 1.435528e-07, 0.00011367941, -6.39699e-05, 8.314424e-07, 1.3839286e-07, 8.17851e-05, -6.359425e-05, 9.439666e-07, 1.3313739e-07, 5.009813e-05, -6.314083e-05, 1.0535388e-06, 1.2779448e-07, 1.8656958e-05, -6.261131e-05, 1.1600637e-06, 1.2237226e-07, -1.2500786e-05, -6.200742e-05, 1.263451e-06, 1.1687877e-07, -4.3338365e-05, -6.133095e-05, 1.3636162e-06, 1.1132208e-07, -7.381995e-05, -6.0583785e-05, 1.4604796e-06, 1.0571017e-07, -0.00010391069, -5.976784e-05, 1.5539671e-06, 1.0005099e-07, -0.00013357666, -5.8885114e-05, 1.6440098e-06, 9.4352416e-08, -0.00016278501, -5.7937654e-05, 1.7305442e-06, 8.8622265e-08, -0.00019150387, -5.6927554e-05, 1.8135123e-06, 8.2868254e-08, -0.00021970247, -5.585697e-05, 1.8928612e-06, 7.7098036e-08, -0.00024735113, -5.4728094e-05, 1.9685433e-06, 7.131915e-08, -0.00027442124, -5.354317e-05, 2.0405166e-06, 6.553904e-08, -0.00030088532, -5.2304473e-05, 2.108744e-06, 5.976505e-08, -0.00032671713, -5.1014315e-05, 2.173194e-06, 5.400438e-08, -0.00035189147, -4.9675047e-05, 2.2338402e-06, 4.8264123e-08, -0.00037638439, -4.828904e-05, 2.2906613e-06, 4.255124e-08, -0.0004001731, -4.68587e-05, 2.343641e-06, 3.687254e-08, -0.00042323608, -4.5386445e-05, 2.3927685e-06, 3.1234695e-08, -0.00044555299, -4.3874727e-05, 2.4380374e-06, 2.5644232e-08, -0.00046710463, -4.2325995e-05, 2.4794467e-06, 2.010751e-08, -0.0004878732, -4.074272e-05, 2.5170002e-06, 1.4630734e-08, -0.00050784205, -3.9127393e-05, 2.5507065e-06, 9.219935e-09, -0.0005269957, -3.7482485e-05, 2.5805787e-06, 3.8809733e-09, -0.00054532, -3.581049e-05, 2.6066346e-06, -1.3804662e-09, -0.0005628021, -3.41139e-05, 2.6288967e-06, -6.5588823e-09, -0.0005794302, -3.239519e-05, 2.6473917e-06, -1.164896e-08, -0.000595194, -3.065684e-05, 2.6621512e-06, -1.6645572e-08, -0.00061008416, -2.8901319e-05, 2.6732105e-06, -2.1543785e-08, -0.0006240928, -2.713108e-05, 2.6806088e-06, -2.6338864e-08, -0.00063721323, -2.5348561e-05, 2.68439e-06, -3.102627e-08, -0.00064943975, -2.3556184e-05, 2.6846017e-06, -3.5601673e-08, -0.0006607681, -2.1756345e-05, 2.6812952e-06, -4.0060936e-08, -0.0006711953, -1.995142e-05, 2.6745254e-06, -4.4400135e-08, -0.0006807191, -1.8143757e-05, 2.6643509e-06, -4.861556e-08, -0.00068933895, -1.6335676e-05, 2.6508335e-06, -5.2703705e-08, -0.0006970551, -1.4529464e-05, 2.634039e-06, -5.666127e-08, -0.0007038691, -1.2727374e-05, 2.6140356e-06, -6.0485185e-08, -0.0007097835, -1.09316225e-05, 2.5908948e-06, -6.417256e-08, -0.0007148021, -9.144388e-06, 2.5646912e-06, -6.772076e-08, -0.0007189297, -7.3678075e-06, 2.535502e-06, -7.112733e-08, -0.0007221721, -5.6039753e-06, 2.503407e-06, -7.439005e-08, -0.00072453613, -3.8549397e-06, 2.4684887e-06, -7.7506904e-08, -0.0007260298, -2.1227038e-06, 2.4308315e-06, -8.047608e-08, -0.00072666194, -4.092206e-07, 2.390523e-06, -8.329599e-08, -0.0007264425, 1.2836073e-06, 2.3476518e-06, -8.5965254e-08, -0.0007253821, 2.9539292e-06, 2.302309e-06, -8.84827e-08, -0.0007234926, 4.5999486e-06, 2.2545876e-06, -9.0847365e-08, -0.0007207865, 6.2199238e-06, 2.2045817e-06, -9.305849e-08, -0.0007172773, 7.81217e-06, 2.1523877e-06, -9.511552e-08, -0.00071297924, 9.375062e-06, 2.0981026e-06, -9.7018095e-08, -0.00070790737, 1.09070315e-05, 2.0418254e-06, -9.876607e-08, -0.0007020776, 1.2406571e-05, 1.9836557e-06, -1.00359486e-07, -0.00069550646, 1.3872235e-05, 1.9236938e-06, -1.0179858e-07, -0.00068821124, 1.5302643e-05, 1.8620416e-06, -1.03083764e-07};
	localparam real hb[0:1199] = {0.011940284, 6.1819783e-06, -8.024018e-06, -8.204753e-09, 0.0119341025, 1.8539538e-05, -8.007101e-06, -2.4590857e-08, 0.011921748, 3.087793e-05, -7.9733045e-06, -4.0907583e-08, 0.01190323, 4.3184416e-05, -7.922693e-06, -5.711045e-08, 0.011878571, 5.5446304e-05, -7.855365e-06, -7.315652e-08, 0.011847793, 6.765098e-05, -7.771447e-06, -8.9004416e-08, 0.01181093, 7.9785925e-05, -7.671095e-06, -1.0461433e-07, 0.011768021, 9.183872e-05, -7.554496e-06, -1.1994803e-07, 0.011719108, 0.00010379708, -7.4218597e-06, -1.349689e-07, 0.011664242, 0.00011564886, -7.273425e-06, -1.4964193e-07, 0.011603478, 0.00012738208, -7.109457e-06, -1.6393372e-07, 0.011536881, 0.00013898496, -6.930243e-06, -1.7781245e-07, 0.011464518, 0.00015044588, -6.7360957e-06, -1.91248e-07, 0.011386461, 0.00016175344, -6.52735e-06, -2.042118e-07, 0.011302792, 0.0001728965, -6.304362e-06, -2.1667695e-07, 0.011213593, 0.00018386412, -6.0675097e-06, -2.2861816e-07, 0.011118958, 0.00019464563, -5.8171895e-06, -2.4001173e-07, 0.01101898, 0.00020523065, -5.5538176e-06, -2.5083557e-07, 0.010913762, 0.00021560903, -5.2778278e-06, -2.6106926e-07, 0.010803408, 0.00022577097, -4.98967e-06, -2.7069387e-07, 0.010688028, 0.00023570693, -4.6898103e-06, -2.7969216e-07, 0.01056774, 0.00024540772, -4.3787304e-06, -2.8804834e-07, 0.010442661, 0.00025486446, -4.0569244e-06, -2.9574826e-07, 0.010312918, 0.0002640686, -3.7248994e-06, -3.027793e-07, 0.010178637, 0.00027301194, -3.383175e-06, -3.0913034e-07, 0.010039951, 0.00028168663, -3.032281e-06, -3.1479172e-07, 0.0098969955, 0.00029008518, -2.672757e-06, -3.1975532e-07, 0.009749913, 0.00029820052, -2.3051512e-06, -3.2401448e-07, 0.009598844, 0.00030602588, -1.93002e-06, -3.2756392e-07, 0.009443936, 0.0003135549, -1.5479261e-06, -3.303998e-07, 0.009285339, 0.00032078158, -1.1594383e-06, -3.325197e-07, 0.009123205, 0.0003277004, -7.6513027e-07, -3.3392251e-07, 0.008957691, 0.00033430613, -3.6557958e-07, -3.3460844e-07, 0.008788953, 0.000340594, 3.863335e-08, -3.3457906e-07, 0.008617151, 0.00034655962, 4.469259e-07, -3.338371e-07, 0.0084424475, 0.00035219904, 8.587143e-07, -3.323867e-07, 0.008265006, 0.00035750863, 1.2734147e-06, -3.3023298e-07, 0.008084994, 0.00036248527, 1.6904436e-06, -3.2738242e-07, 0.0079025775, 0.0003671262, 2.1092192e-06, -3.2384258e-07, 0.007717924, 0.00037142902, 2.529162e-06, -3.1962207e-07, 0.0075312047, 0.00037539183, 2.9496955e-06, -3.1473067e-07, 0.007342589, 0.0003790131, 3.3702477e-06, -3.0917906e-07, 0.0071522486, 0.00038229168, 3.7902503e-06, -3.0297903e-07, 0.0069603547, 0.00038522683, 4.2091415e-06, -2.9614327e-07, 0.0067670792, 0.0003878182, 4.626366e-06, -2.886854e-07, 0.006572594, 0.00039006592, 5.0413737e-06, -2.8061996e-07, 0.0063770707, 0.0003919704, 5.4536245e-06, -2.7196222e-07, 0.006180681, 0.0003935325, 5.8625856e-06, -2.6272835e-07, 0.005983595, 0.00039475344, 6.267733e-06, -2.529353e-07, 0.0057859835, 0.00039563482, 6.668553e-06, -2.4260066e-07, 0.0055880165, 0.00039617866, 7.0645415e-06, -2.3174275e-07, 0.005389861, 0.00039638727, 7.4552063e-06, -2.2038053e-07, 0.0051916847, 0.0003962634, 7.840066e-06, -2.0853356e-07, 0.0049936525, 0.0003958101, 8.218651e-06, -1.9622199e-07, 0.004795929, 0.00039503071, 8.590505e-06, -1.8346643e-07, 0.0045986753, 0.00039392908, 8.955183e-06, -1.7028802e-07, 0.0044020526, 0.00039250925, 9.312257e-06, -1.5670835e-07, 0.0042062183, 0.00039077562, 9.6613085e-06, -1.4274937e-07, 0.004011329, 0.0003887329, 1.0001936e-05, -1.2843343e-07, 0.0038175362, 0.00038638615, 1.0333753e-05, -1.1378318e-07, 0.0036249922, 0.00038374067, 1.0656387e-05, -9.882157e-08, 0.0034338445, 0.00038080206, 1.096948e-05, -8.3571805e-08, 0.003244238, 0.0003775762, 1.1272693e-05, -6.805727e-08, 0.0030563152, 0.00037406923, 1.15656985e-05, -5.2301523e-08, 0.0028702146, 0.00037028757, 1.1848189e-05, -3.6328274e-08, 0.0026860721, 0.00036623792, 1.2119873e-05, -2.016131e-08, 0.0025040202, 0.0003619271, 1.2380473e-05, -3.8244825e-09, 0.0023241874, 0.00035736224, 1.2629732e-05, 1.265834e-08, 0.0021466992, 0.0003525507, 1.2867406e-05, 2.92633e-08, 0.0019716767, 0.00034749997, 1.3093272e-05, 4.5966587e-08, 0.0017992377, 0.00034221783, 1.33071235e-05, 6.274448e-08, 0.0016294961, 0.0003367121, 1.35087685e-05, 7.957337e-08, 0.0014625615, 0.00033099094, 1.3698036e-05, 9.6429794e-08, 0.0012985397, 0.00032506252, 1.387477e-05, 1.13290476e-07, 0.0011375322, 0.00031893523, 1.4038833e-05, 1.3013234e-07, 0.0009796362, 0.00031261757, 1.4190105e-05, 1.4693258e-07, 0.0008249449, 0.0003061182, 1.43284815e-05, 1.6366863e-07, 0.00067354686, 0.00029944582, 1.4453879e-05, 1.8031824e-07, 0.0005255264, 0.00029260933, 1.4566228e-05, 1.9685949e-07, 0.0003809634, 0.0002856176, 1.46654775e-05, 2.1327081e-07, 0.00023993319, 0.00027847965, 1.4751593e-05, 2.2953101e-07, 0.00010250661, 0.00027120457, 1.4824558e-05, 2.4561933e-07, -3.1250034e-05, 0.00026380146, 1.488437e-05, 2.615154e-07, -0.00016127502, 0.00025627948, 1.4931046e-05, 2.7719932e-07, -0.00028751124, 0.00024864782, 1.4964618e-05, 2.926517e-07, -0.0004099061, 0.00024091572, 1.4985132e-05, 3.0785355e-07, -0.0005284117, 0.00023309235, 1.49926545e-05, 3.2278655e-07, -0.00064298476, 0.00022518694, 1.4987263e-05, 3.374328e-07, -0.00075358653, 0.00021720871, 1.4969053e-05, 3.5177496e-07, -0.00086018286, 0.00020916681, 1.4938134e-05, 3.6579627e-07, -0.00096274423, 0.00020107039, 1.4894629e-05, 3.794806e-07, -0.0010612457, 0.00019292852, 1.4838679e-05, 3.9281244e-07, -0.0011556667, 0.00018475026, 1.4770433e-05, 4.0577677e-07, -0.0012459913, 0.00017654453, 1.469006e-05, 4.183593e-07, -0.0013322082, 0.00016832027, 1.4597737e-05, 4.3054638e-07, -0.00141431, 0.00016008626, 1.4493659e-05, 4.42325e-07, -0.0014922943, 0.0001518512, 1.4378028e-05, 4.5368273e-07, -0.0015661624, 0.0001436237, 1.4251062e-05, 4.6460795e-07, -0.0016359206, 0.00013541225, 1.41129885e-05, 4.7508965e-07, -0.0017015787, 0.00012722521, 1.3964048e-05, 4.851175e-07, -0.0017631513, 0.00011907082, 1.3804491e-05, 4.946818e-07, -0.0018206564, 0.00011095717, 1.3634577e-05, 5.0377366e-07, -0.0018741165, 0.00010289221, 1.3454577e-05, 5.123848e-07, -0.001923558, 9.488373e-05, 1.3264772e-05, 5.205078e-07, -0.001969011, 8.693937e-05, 1.306545e-05, 5.281357e-07, -0.0020105094, 7.906658e-05, 1.2856909e-05, 5.352623e-07, -0.0020480906, 7.1272654e-05, 1.2639454e-05, 5.4188234e-07, -0.0020817963, 6.3564694e-05, 1.2413399e-05, 5.4799096e-07, -0.0021116708, 5.594962e-05, 1.2179065e-05, 5.535842e-07, -0.0021377625, 4.8434144e-05, 1.1936777e-05, 5.5865866e-07, -0.0021601226, 4.1024792e-05, 1.1686869e-05, 5.6321176e-07, -0.002178806, 3.3727883e-05, 1.1429678e-05, 5.6724144e-07, -0.0021938703, 2.654952e-05, 1.116555e-05, 5.707466e-07, -0.0022053763, 1.94956e-05, 1.08948325e-05, 5.737265e-07, -0.0022133875, 1.257179e-05, 1.0617877e-05, 5.761812e-07, -0.0022179708, 5.7835446e-06, 1.033504e-05, 5.781115e-07, -0.0022191945, -8.6391225e-07, 1.0046682e-05, 5.795188e-07, -0.002217131, -7.365586e-06, 9.753164e-06, 5.8040507e-07, -0.002211854, -1.3716714e-05, 9.45485e-06, 5.80773e-07, -0.0022034403, -1.991277e-05, 9.152107e-06, 5.806259e-07, -0.0021919678, -2.5949465e-05, 8.845302e-06, 5.799676e-07, -0.0021775179, -3.1822747e-05, 8.534802e-06, 5.7880266e-07, -0.002160173, -3.7528807e-05, 8.220977e-06, 5.7713606e-07, -0.0021400177, -4.3064083e-05, 7.904194e-06, 5.7497346e-07, -0.002117138, -4.8425245e-05, 7.58482e-06, 5.7232114e-07, -0.002091622, -5.3609227e-05, 7.263224e-06, 5.691858e-07, -0.0020635587, -5.8613183e-05, 6.9397693e-06, 5.655747e-07, -0.0020330392, -6.3434534e-05, 6.6148195e-06, 5.614956e-07, -0.002000155, -6.8070935e-05, 6.288736e-06, 5.569569e-07, -0.0019649994, -7.2520284e-05, 5.961877e-06, 5.5196716e-07, -0.0019276662, -7.678073e-05, 5.634597e-06, 5.4653583e-07, -0.0018882505, -8.085066e-05, 5.3072476e-06, 5.406724e-07, -0.0018468476, -8.472871e-05, 4.980177e-06, 5.34387e-07, -0.0018035539, -8.841373e-05, 4.6537284e-06, 5.2769025e-07, -0.0017584661, -9.190485e-05, 4.32824e-06, 5.2059295e-07, -0.0017116815, -9.5201394e-05, 4.0040454e-06, 5.131064e-07, -0.0016632973, -9.830295e-05, 3.681473e-06, 5.0524216e-07, -0.001613411, -0.00010120933, 3.360845e-06, 4.970123e-07, -0.0015621204, -0.00010392056, 3.0424783e-06, 4.88429e-07, -0.001509523, -0.0001064369, 2.7266829e-06, 4.79505e-07, -0.001455716, -0.00010875883, 2.413762e-06, 4.7025296e-07, -0.0014007965, -0.00011088706, 2.1040125e-06, 4.6068612e-07, -0.001344861, -0.0001128225, 1.7977234e-06, 4.508178e-07, -0.0012880058, -0.00011456626, 1.4951765e-06, 4.4066155e-07, -0.0012303265, -0.00011611969, 1.1966463e-06, 4.302312e-07, -0.0011719177, -0.00011748432, 9.023985e-07, 4.1954067e-07, -0.0011128733, -0.00011866187, 6.126912e-07, 4.0860408e-07, -0.0010532866, -0.000119654265, 3.2777407e-07, 3.9743568e-07, -0.0009932496, -0.000120463614, 4.7888012e-08, 3.8604986e-07, -0.00093285315, -0.0001210922, -2.2673481e-07, 3.7446114e-07, -0.0008721871, -0.00012154251, -4.958712e-07, 3.62684e-07, -0.00081133994, -0.00012181716, -7.5930694e-07, 3.5073316e-07, -0.0007503987, -0.00012191897, -1.0168372e-06, 3.386232e-07, -0.00068944925, -0.000121850906, -1.2682666e-06, 3.2636893e-07, -0.0006285756, -0.00012161609, -1.5134091e-06, 3.1398497e-07, -0.00056786044, -0.00012121779, -1.7520883e-06, 3.0148607e-07, -0.00050738454, -0.00012065941, -1.9841377e-06, 2.8888687e-07, -0.0004472271, -0.00011994451, -2.2094002e-06, 2.7620203e-07, -0.0003874655, -0.00011907677, -2.427729e-06, 2.6344605e-07, -0.00032817517, -0.000118059994, -2.6389869e-06, 2.506335e-07, -0.0002694297, -0.0001168981, -2.8430466e-06, 2.3777866e-07, -0.00021130059, -0.00011559514, -3.039791e-06, 2.2489587e-07, -0.00015385737, -0.00011415523, -3.2291125e-06, 2.1199925e-07, -9.7167474e-05, -0.000112582624, -3.4109146e-06, 1.9910277e-07, -4.129615e-05, -0.00011088165, -3.5851092e-06, 1.8622028e-07, 1.3693514e-05, -0.000109056724, -3.7516195e-06, 1.7336544e-07, 6.7740664e-05, -0.000107112355, -3.910378e-06, 1.6055168e-07, 0.00012078672, -0.0001050531, -4.0613268e-06, 1.4779228e-07, 0.00017277538, -0.0001028836, -4.2044185e-06, 1.3510027e-07, 0.00022365272, -0.00010060855, -4.3396144e-06, 1.2248844e-07, 0.00027336713, -9.823271e-05, -4.4668873e-06, 1.09969385e-07, 0.00032186942, -9.576087e-05, -4.5862175e-06, 9.755537e-08, 0.00036911282, -9.319787e-05, -4.6975956e-06, 8.525845e-08, 0.00041505293, -9.054859e-05, -4.8010224e-06, 7.309037e-08, 0.00045964782, -8.781791e-05, -4.896506e-06, 6.106258e-08, 0.0005028581, -8.501077e-05, -4.984066e-06, 4.9186248e-08, 0.0005446467, -8.21321e-05, -5.063729e-06, 3.7472216e-08, 0.0005849791, -7.9186844e-05, -5.1355314e-06, 2.593101e-08, 0.00062382326, -7.617996e-05, -5.199517e-06, 1.45728265e-08, 0.0006611496, -7.311639e-05, -5.2557402e-06, 3.4075192e-09, 0.00069693103, -7.000107e-05, -5.3042622e-06, -7.5554e-09, 0.0007311429, -6.683892e-05, -5.3451527e-06, -1.8306773e-08, 0.0007637629, -6.363485e-05, -5.3784884e-06, -2.8837803e-08, 0.00079477153, -6.039373e-05, -5.4043558e-06, -3.914006e-08, 0.0008241513, -5.712041e-05, -5.422847e-06, -4.920548e-08, 0.0008518874, -5.3819695e-05, -5.4340626e-06, -5.902638e-08, 0.0008779672, -5.0496346e-05, -5.4381094e-06, -6.859546e-08, 0.00090238074, -4.715509e-05, -5.4351017e-06, -7.79058e-08, 0.0009251201, -4.3800588e-05, -5.4251605e-06, -8.6950884e-08, 0.00094617985, -4.0437444e-05, -5.408412e-06, -9.572456e-08, 0.0009655569, -3.7070215e-05, -5.384991e-06, -1.0422109e-07, 0.0009832501, -3.3703367e-05, -5.3550352e-06, -1.1243513e-07, 0.000999261, -3.034132e-05, -5.3186905e-06, -1.2036173e-07, 0.001013593, -2.6988402e-05, -5.276107e-06, -1.2799634e-07, 0.0010262517, -2.3648865e-05, -5.22744e-06, -1.3533482e-07, 0.0010372448, -2.032688e-05, -5.17285e-06, -1.423734e-07, 0.0010465821, -1.7026527e-05, -5.112502e-06, -1.4910871e-07, 0.0010542755, -1.3751798e-05, -5.046566e-06, -1.5553783e-07, 0.0010603388, -1.050659e-05, -4.9752152e-06, -1.6165818e-07, 0.0010647877, -7.2947e-06, -4.898627e-06, -1.6746759e-07, 0.0010676397, -4.119824e-06, -4.8169827e-06, -1.7296428e-07, 0.0010689143, -9.855555e-07, -4.730466e-06, -1.7814686e-07, 0.0010686326, 2.1046212e-06, -4.639265e-06, -1.8301432e-07, 0.0010668176, 5.147331e-06, -4.5435704e-06, -1.8756604e-07, 0.0010634938, 8.139311e-06, -4.4435737e-06, -1.9180179e-07, 0.0010586872, 1.1077412e-05, -4.3394707e-06, -1.9572165e-07, 0.0010524258, 1.3958604e-05, -4.2314587e-06, -1.9932614e-07, 0.0010447387, 1.6779974e-05, -4.119736e-06, -2.026161e-07, 0.0010356563, 1.953873e-05, -4.0045024e-06, -2.0559277e-07, 0.0010252108, 2.2232203e-05, -3.8859603e-06, -2.0825766e-07, 0.0010134354, 2.4857845e-05, -3.7643117e-06, -2.1061268e-07, 0.0010003647, 2.741324e-05, -3.6397594e-06, -2.1266008e-07, 0.0009860343, 2.989609e-05, -3.512507e-06, -2.1440243e-07, 0.000970481, 3.230423e-05, -3.3827585e-06, -2.1584259e-07, 0.0009537428, 3.4635617e-05, -3.2507169e-06, -2.1698379e-07, 0.0009358585, 3.6888345e-05, -3.116586e-06, -2.1782952e-07, 0.00091686787, 3.906063e-05, -2.9805683e-06, -2.1838359e-07, 0.00089681154, 4.1150815e-05, -2.842866e-06, -2.1865007e-07, 0.000875731, 4.3157386e-05, -2.7036797e-06, -2.1863337e-07, 0.0008536683, 4.5078945e-05, -2.5632094e-06, -2.1833812e-07, 0.00083066645, 4.691423e-05, -2.421653e-06, -2.177692e-07, 0.00080676866, 4.86621e-05, -2.2792071e-06, -2.1693181e-07, 0.00078201905, 5.0321552e-05, -2.1360665e-06, -2.1583132e-07, 0.000756462, 5.1891704e-05, -1.9924237e-06, -2.1447337e-07, 0.00073014235, 5.337181e-05, -1.8484684e-06, -2.1286382e-07, 0.0007031053, 5.4761233e-05, -1.7043886e-06, -2.1100877e-07, 0.00067539635, 5.6059478e-05, -1.5603694e-06, -2.0891444e-07, 0.0006470611, 5.7266167e-05, -1.4165925e-06, -2.0658733e-07, 0.00061814545, 5.8381043e-05, -1.273237e-06, -2.0403407e-07, 0.0005886954, 5.940397e-05, -1.1304786e-06, -2.012615e-07, 0.0005587568, 6.0334933e-05, -9.884898e-07, -1.9827658e-07, 0.0005283758, 6.117403e-05, -8.474391e-07, -1.9508646e-07, 0.0004975981, 6.192149e-05, -7.074916e-07, -1.9169838e-07, 0.0004664695, 6.257763e-05, -5.6880845e-07, -1.8811977e-07, 0.0004350356, 6.31429e-05, -4.3154677e-07, -1.8435814e-07, 0.00040334166, 6.3617845e-05, -2.958595e-07, -1.8042111e-07, 0.0003714327, 6.400313e-05, -1.6189534e-07, -1.763164e-07, 0.00033935334, 6.4299515e-05, -2.9798583e-08, -1.7205184e-07, 0.00030714786, 6.450787e-05, 1.0029098e-07, -1.6763529e-07, 0.00027485998, 6.4629145e-05, 2.2823818e-07, -1.6307472e-07, 0.00024253305, 6.466442e-05, 3.5391255e-07, -1.5837811e-07, 0.00021020972, 6.461484e-05, 4.7718845e-07, -1.5355353e-07, 0.00017793213, 6.4481654e-05, 5.979451e-07, -1.4860906e-07, 0.00014574177, 6.42662e-05, 7.1606667e-07, -1.435528e-07, 0.00011367941, 6.39699e-05, 8.314424e-07, -1.3839286e-07, 8.17851e-05, 6.359425e-05, 9.439666e-07, -1.3313739e-07, 5.009813e-05, 6.314083e-05, 1.0535388e-06, -1.2779448e-07, 1.8656958e-05, 6.261131e-05, 1.1600637e-06, -1.2237226e-07, -1.2500786e-05, 6.200742e-05, 1.263451e-06, -1.1687877e-07, -4.3338365e-05, 6.133095e-05, 1.3636162e-06, -1.1132208e-07, -7.381995e-05, 6.0583785e-05, 1.4604796e-06, -1.0571017e-07, -0.00010391069, 5.976784e-05, 1.5539671e-06, -1.0005099e-07, -0.00013357666, 5.8885114e-05, 1.6440098e-06, -9.4352416e-08, -0.00016278501, 5.7937654e-05, 1.7305442e-06, -8.8622265e-08, -0.00019150387, 5.6927554e-05, 1.8135123e-06, -8.2868254e-08, -0.00021970247, 5.585697e-05, 1.8928612e-06, -7.7098036e-08, -0.00024735113, 5.4728094e-05, 1.9685433e-06, -7.131915e-08, -0.00027442124, 5.354317e-05, 2.0405166e-06, -6.553904e-08, -0.00030088532, 5.2304473e-05, 2.108744e-06, -5.976505e-08, -0.00032671713, 5.1014315e-05, 2.173194e-06, -5.400438e-08, -0.00035189147, 4.9675047e-05, 2.2338402e-06, -4.8264123e-08, -0.00037638439, 4.828904e-05, 2.2906613e-06, -4.255124e-08, -0.0004001731, 4.68587e-05, 2.343641e-06, -3.687254e-08, -0.00042323608, 4.5386445e-05, 2.3927685e-06, -3.1234695e-08, -0.00044555299, 4.3874727e-05, 2.4380374e-06, -2.5644232e-08, -0.00046710463, 4.2325995e-05, 2.4794467e-06, -2.010751e-08, -0.0004878732, 4.074272e-05, 2.5170002e-06, -1.4630734e-08, -0.00050784205, 3.9127393e-05, 2.5507065e-06, -9.219935e-09, -0.0005269957, 3.7482485e-05, 2.5805787e-06, -3.8809733e-09, -0.00054532, 3.581049e-05, 2.6066346e-06, 1.3804662e-09, -0.0005628021, 3.41139e-05, 2.6288967e-06, 6.5588823e-09, -0.0005794302, 3.239519e-05, 2.6473917e-06, 1.164896e-08, -0.000595194, 3.065684e-05, 2.6621512e-06, 1.6645572e-08, -0.00061008416, 2.8901319e-05, 2.6732105e-06, 2.1543785e-08, -0.0006240928, 2.713108e-05, 2.6806088e-06, 2.6338864e-08, -0.00063721323, 2.5348561e-05, 2.68439e-06, 3.102627e-08, -0.00064943975, 2.3556184e-05, 2.6846017e-06, 3.5601673e-08, -0.0006607681, 2.1756345e-05, 2.6812952e-06, 4.0060936e-08, -0.0006711953, 1.995142e-05, 2.6745254e-06, 4.4400135e-08, -0.0006807191, 1.8143757e-05, 2.6643509e-06, 4.861556e-08, -0.00068933895, 1.6335676e-05, 2.6508335e-06, 5.2703705e-08, -0.0006970551, 1.4529464e-05, 2.634039e-06, 5.666127e-08, -0.0007038691, 1.2727374e-05, 2.6140356e-06, 6.0485185e-08, -0.0007097835, 1.09316225e-05, 2.5908948e-06, 6.417256e-08, -0.0007148021, 9.144388e-06, 2.5646912e-06, 6.772076e-08, -0.0007189297, 7.3678075e-06, 2.535502e-06, 7.112733e-08, -0.0007221721, 5.6039753e-06, 2.503407e-06, 7.439005e-08, -0.00072453613, 3.8549397e-06, 2.4684887e-06, 7.7506904e-08, -0.0007260298, 2.1227038e-06, 2.4308315e-06, 8.047608e-08, -0.00072666194, 4.092206e-07, 2.390523e-06, 8.329599e-08, -0.0007264425, -1.2836073e-06, 2.3476518e-06, 8.5965254e-08, -0.0007253821, -2.9539292e-06, 2.302309e-06, 8.84827e-08, -0.0007234926, -4.5999486e-06, 2.2545876e-06, 9.0847365e-08, -0.0007207865, -6.2199238e-06, 2.2045817e-06, 9.305849e-08, -0.0007172773, -7.81217e-06, 2.1523877e-06, 9.511552e-08, -0.00071297924, -9.375062e-06, 2.0981026e-06, 9.7018095e-08, -0.00070790737, -1.09070315e-05, 2.0418254e-06, 9.876607e-08, -0.0007020776, -1.2406571e-05, 1.9836557e-06, 1.00359486e-07, -0.00069550646, -1.3872235e-05, 1.9236938e-06, 1.0179858e-07, -0.00068821124, -1.5302643e-05, 1.8620416e-06, 1.03083764e-07};
endpackage
`endif
