`ifndef COEFFICIENTS_FX_SV_
`define COEFFICIENTS_FX_SV_
package Coefficients_Fx;
	localparam N = 3;
	localparam M = 3;
	localparam COEFF_BIAS = 48;
	localparam logic signed[63:0] Lfr[0:2] = {64'd261058313901802, 64'd269039775171046, 64'd269039775171046};
	localparam logic signed[63:0] Lfi[0:2] = {64'd0, 64'd30680189886302, - 64'd30680189886302};
	localparam logic signed[63:0] Lbr[0:2] = {64'd261058313901802, 64'd269039775171046, 64'd269039775171046};
	localparam logic signed[63:0] Lbi[0:2] = {64'd0, 64'd30680189886302, - 64'd30680189886302};
	localparam logic signed[63:0] Wfr[0:2] = {- 64'd686598368623, 64'd433640635081, 64'd433640635081};
	localparam logic signed[63:0] Wfi[0:2] = {64'd0, - 64'd811113628749, 64'd811113628749};
	localparam logic signed[63:0] Wbr[0:2] = {64'd686598368623, - 64'd433640635081, - 64'd433640635081};
	localparam logic signed[63:0] Wbi[0:2] = {64'd0, 64'd811113628749, - 64'd811113628749};
	localparam logic signed[63:0] Ffr[0:2][0:74] = '{
		'{- 64'd2302183503407588, 64'd345904573056852, - 64'd94577992473653, - 64'd2135195642310809, 64'd320814538004102, - 64'd87717819665262, - 64'd1980320171782550, 64'd297544397534951, - 64'd81355246454094, - 64'd1836678524935849, 64'd275962146401561, - 64'd75454179673682, - 64'd1703455861343890, 64'd255945354298297, - 64'd69981144159410, - 64'd1579896444669438, 64'd237380471347538, - 64'd64905092852906, - 64'd1465299355575864, 64'd220162183961760, - 64'd60197230680428, - 64'd1359014515600282, 64'd204192817427879, - 64'd55830851206161, - 64'd1260438999433276, 64'd189381781824880, - 64'd51781185133787, - 64'd1169013614685802, 64'd175645058131558, - 64'd48025259796928, - 64'd1084219729741160, 64'd162904721609211, - 64'd44541768841391, - 64'd1005576331697337, 64'd151088499755556, - 64'd41310951359952, - 64'd932637297710195, 64'd140129362322264, - 64'd38314479794040, - 64'd864988864258566, 64'd129965141070389, - 64'd35535355966434, - 64'd802247279975093, 64'd120538177106673, - 64'd32957814655168, - 64'd744056628727935, 64'd111794993800149, - 64'd30567234161674, - 64'd690086810604292, 64'd103685993423601, - 64'd28350053365813, - 64'd640031669342381, 64'd96165175798997, - 64'd26293694797294, - 64'd593607255589311, 64'd89189877350849, - 64'd24386493287061, - 64'd550550216132783, 64'd82720529087230, - 64'd22617629793934, - 64'd510616299969148, 64'd76720432135521, - 64'd20977070031092, - 64'd473578972733160, 64'd71155549559580, - 64'd19455507544269, - 64'd439228131629457, 64'd65994313277358, - 64'd18044310918734, - 64'd407368913575912, 64'd61207444983660, - 64'd16735474815607, - 64'd377820589797780, 64'd56767790062194, - 64'd15521574559714},
		'{64'd1194733174907733, - 64'd196745053762742, - 64'd19558774927113, 64'd1091854361667905, - 64'd213796329652344, - 64'd12910391622595, 64'd981539738675941, - 64'd226619560737254, - 64'd6578899337396, 64'd865869366263096, - 64'd235352467665655, - 64'd628260878998, 64'd746842370399115, - 64'd240179086059323, 64'd4887595867794, 64'd626355321810053, - 64'd241323769247672, 64'd9924776034165, 64'd506183644970437, - 64'd239045080261807, 64'd14449277222949, 64'd387966088324595, - 64'd233629665829313, 64'd18436722602651, 64'd273192242411343, - 64'd225386198447957, 64'd21871980748900, 64'd163193051399847, - 64'd214639465259820, 64'd24748685931934, 64'd59134226199680, - 64'd201724674550048, 64'd27068672904946, - 64'd37987565983178, - 64'd186982042405970, 64'd28841340383285, - 64'd127345889852109, - 64'd170751713536614, 64'd30082957333395, - 64'd208283286974387, - 64'd153369061606049, 64'd30815925929228, - 64'd280307776928200, - 64'd135160405804480, 64'd31068014600502, - 64'd343087330259404, - 64'd116439171886633, 64'd30871574010424, - 64'd396442540850866, - 64'd97502517655162, 64'd30262748079906, - 64'd440337733251421, - 64'd78628434953589, 64'd29280691340780, - 64'd474870744605419, - 64'd60073332742995, 64'd27966802972162, - 64'd500261621297886, - 64'd42070098841254, 64'd26363986871690, - 64'd516840467547726, - 64'd24826631463055, 64'd24515946056310, - 64'd525034677232123, - 64'd8524825860936, 64'd22466518594256, - 64'd525355771520235, 64'd6680003832020, 64'd20259061158714, - 64'd518386053759184, 64'd20659291994046, 64'd17935885181011, - 64'd504765279825352, 64'd33311006438020, 64'd15537749482665},
		'{64'd1194733174907733, - 64'd196745053762742, - 64'd19558774927113, 64'd1091854361667905, - 64'd213796329652344, - 64'd12910391622595, 64'd981539738675941, - 64'd226619560737254, - 64'd6578899337396, 64'd865869366263096, - 64'd235352467665655, - 64'd628260878998, 64'd746842370399115, - 64'd240179086059323, 64'd4887595867794, 64'd626355321810053, - 64'd241323769247672, 64'd9924776034165, 64'd506183644970437, - 64'd239045080261808, 64'd14449277222949, 64'd387966088324595, - 64'd233629665829313, 64'd18436722602651, 64'd273192242411343, - 64'd225386198447957, 64'd21871980748900, 64'd163193051399847, - 64'd214639465259820, 64'd24748685931934, 64'd59134226199680, - 64'd201724674550048, 64'd27068672904946, - 64'd37987565983178, - 64'd186982042405970, 64'd28841340383285, - 64'd127345889852109, - 64'd170751713536614, 64'd30082957333395, - 64'd208283286974387, - 64'd153369061606049, 64'd30815925929228, - 64'd280307776928200, - 64'd135160405804480, 64'd31068014600502, - 64'd343087330259404, - 64'd116439171886633, 64'd30871574010424, - 64'd396442540850866, - 64'd97502517655162, 64'd30262748079906, - 64'd440337733251421, - 64'd78628434953589, 64'd29280691340780, - 64'd474870744605419, - 64'd60073332742995, 64'd27966802972162, - 64'd500261621297886, - 64'd42070098841254, 64'd26363986871690, - 64'd516840467547726, - 64'd24826631463055, 64'd24515946056310, - 64'd525034677232123, - 64'd8524825860936, 64'd22466518594256, - 64'd525355771520235, 64'd6680003832020, 64'd20259061158714, - 64'd518386053759184, 64'd20659291994046, 64'd17935885181011, - 64'd504765279825352, 64'd33311006438020, 64'd15537749482665}};
	localparam logic signed[63:0] Ffi[0:2][0:74] = '{
		'{64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0},
		'{64'd459614617670948, 64'd236180802864224, - 64'd53067997093561, 64'd569532879783993, 64'd204301835870795, - 64'd52855387393211, 64'd663381517092044, 64'd171972686754111, - 64'd51927510495402, 64'd741059977026027, 64'd139674092112747, - 64'd50350506447889, 64'd802698871570680, 64'd107850538956602, - 64'd48194565130026, 64'd848640943034727, 64'd76906817930726, - 64'd45532653550627, 64'd879420514097390, 64'd47205382502847, - 64'd42439299579991, 64'd895741819343958, 64'd19064490578595, - 64'd38989444734119, 64'd898456601372454, - 64'd7242904060338, - 64'd35257376733643, 64'd888541336176843, - 64'd31489551041779, - 64'd31315750657421, 64'd867074430460488, - 64'd53493640748254, - 64'd27234705627979, 64'd835213708385532, - 64'd73117932686057, - 64'd23081082127544, 64'd794174477598151, - 64'd90268332318900, - 64'd18917743271502, 64'd745208434756558, - 64'd104891977155066, - 64'd14803001680187, 64'd689583639782946, - 64'd116974895134814, - 64'd10790152006959, 64'd628565756194885, - 64'd126539299582327, - 64'd6927107714744, 64'd563400722650966, - 64'd133640585224329, - 64'd3256139356123, 64'd495298988741795, - 64'd138364089105400, 64'd186289587403, 64'd425421416506145, - 64'd140821678725097, 64'd3369594306864, 64'd354866918548485, - 64'd141148227467154, 64'd6269053615551, 64'd284661874330815, - 64'd139498034473248, 64'd8865714912952, 64'd215751338517271, - 64'd136041242623042, 64'd11146226438403, 64'd148992029427446, - 64'd130960304309206, 64'd13102604553515, 64'd85147061921491, - 64'd124446540332005, 64'd14731944114389, 64'd24882367569355, - 64'd116696832572115, 64'd16036080181081},
		'{- 64'd459614617670948, - 64'd236180802864224, 64'd53067997093561, - 64'd569532879783993, - 64'd204301835870795, 64'd52855387393211, - 64'd663381517092044, - 64'd171972686754111, 64'd51927510495402, - 64'd741059977026027, - 64'd139674092112747, 64'd50350506447889, - 64'd802698871570680, - 64'd107850538956602, 64'd48194565130026, - 64'd848640943034728, - 64'd76906817930726, 64'd45532653550627, - 64'd879420514097390, - 64'd47205382502847, 64'd42439299579991, - 64'd895741819343958, - 64'd19064490578595, 64'd38989444734119, - 64'd898456601372454, 64'd7242904060338, 64'd35257376733643, - 64'd888541336176843, 64'd31489551041779, 64'd31315750657421, - 64'd867074430460488, 64'd53493640748254, 64'd27234705627979, - 64'd835213708385532, 64'd73117932686057, 64'd23081082127544, - 64'd794174477598151, 64'd90268332318900, 64'd18917743271502, - 64'd745208434756558, 64'd104891977155066, 64'd14803001680187, - 64'd689583639782946, 64'd116974895134814, 64'd10790152006959, - 64'd628565756194885, 64'd126539299582327, 64'd6927107714744, - 64'd563400722650966, 64'd133640585224329, 64'd3256139356123, - 64'd495298988741795, 64'd138364089105400, - 64'd186289587403, - 64'd425421416506145, 64'd140821678725097, - 64'd3369594306864, - 64'd354866918548485, 64'd141148227467154, - 64'd6269053615551, - 64'd284661874330815, 64'd139498034473249, - 64'd8865714912952, - 64'd215751338517271, 64'd136041242623042, - 64'd11146226438403, - 64'd148992029427446, 64'd130960304309206, - 64'd13102604553515, - 64'd85147061921491, 64'd124446540332005, - 64'd14731944114389, - 64'd24882367569355, 64'd116696832572115, - 64'd16036080181081}};
	localparam logic signed[63:0] Fbr[0:2][0:74] = '{
		'{64'd2302183503407588, 64'd345904573056852, 64'd94577992473653, 64'd2135195642310809, 64'd320814538004102, 64'd87717819665262, 64'd1980320171782550, 64'd297544397534951, 64'd81355246454094, 64'd1836678524935849, 64'd275962146401561, 64'd75454179673682, 64'd1703455861343890, 64'd255945354298297, 64'd69981144159410, 64'd1579896444669438, 64'd237380471347538, 64'd64905092852906, 64'd1465299355575864, 64'd220162183961760, 64'd60197230680428, 64'd1359014515600282, 64'd204192817427879, 64'd55830851206161, 64'd1260438999433276, 64'd189381781824880, 64'd51781185133787, 64'd1169013614685802, 64'd175645058131558, 64'd48025259796928, 64'd1084219729741160, 64'd162904721609211, 64'd44541768841391, 64'd1005576331697337, 64'd151088499755556, 64'd41310951359952, 64'd932637297710195, 64'd140129362322264, 64'd38314479794040, 64'd864988864258566, 64'd129965141070389, 64'd35535355966434, 64'd802247279975093, 64'd120538177106673, 64'd32957814655168, 64'd744056628727935, 64'd111794993800149, 64'd30567234161674, 64'd690086810604292, 64'd103685993423601, 64'd28350053365813, 64'd640031669342381, 64'd96165175798997, 64'd26293694797294, 64'd593607255589311, 64'd89189877350849, 64'd24386493287061, 64'd550550216132783, 64'd82720529087230, 64'd22617629793934, 64'd510616299969148, 64'd76720432135521, 64'd20977070031092, 64'd473578972733160, 64'd71155549559580, 64'd19455507544269, 64'd439228131629457, 64'd65994313277358, 64'd18044310918734, 64'd407368913575912, 64'd61207444983660, 64'd16735474815607, 64'd377820589797780, 64'd56767790062194, 64'd15521574559714},
		'{- 64'd1194733174907733, - 64'd196745053762742, 64'd19558774927113, - 64'd1091854361667905, - 64'd213796329652344, 64'd12910391622595, - 64'd981539738675941, - 64'd226619560737254, 64'd6578899337396, - 64'd865869366263096, - 64'd235352467665655, 64'd628260878998, - 64'd746842370399115, - 64'd240179086059323, - 64'd4887595867794, - 64'd626355321810053, - 64'd241323769247672, - 64'd9924776034165, - 64'd506183644970437, - 64'd239045080261807, - 64'd14449277222949, - 64'd387966088324595, - 64'd233629665829313, - 64'd18436722602651, - 64'd273192242411343, - 64'd225386198447957, - 64'd21871980748900, - 64'd163193051399847, - 64'd214639465259820, - 64'd24748685931934, - 64'd59134226199680, - 64'd201724674550048, - 64'd27068672904946, 64'd37987565983178, - 64'd186982042405970, - 64'd28841340383285, 64'd127345889852109, - 64'd170751713536614, - 64'd30082957333395, 64'd208283286974387, - 64'd153369061606049, - 64'd30815925929228, 64'd280307776928200, - 64'd135160405804480, - 64'd31068014600502, 64'd343087330259404, - 64'd116439171886633, - 64'd30871574010424, 64'd396442540850866, - 64'd97502517655162, - 64'd30262748079906, 64'd440337733251421, - 64'd78628434953589, - 64'd29280691340780, 64'd474870744605419, - 64'd60073332742995, - 64'd27966802972162, 64'd500261621297886, - 64'd42070098841254, - 64'd26363986871690, 64'd516840467547726, - 64'd24826631463055, - 64'd24515946056310, 64'd525034677232123, - 64'd8524825860936, - 64'd22466518594256, 64'd525355771520235, 64'd6680003832020, - 64'd20259061158714, 64'd518386053759184, 64'd20659291994046, - 64'd17935885181011, 64'd504765279825352, 64'd33311006438020, - 64'd15537749482665},
		'{- 64'd1194733174907733, - 64'd196745053762742, 64'd19558774927113, - 64'd1091854361667905, - 64'd213796329652344, 64'd12910391622595, - 64'd981539738675941, - 64'd226619560737254, 64'd6578899337396, - 64'd865869366263096, - 64'd235352467665655, 64'd628260878998, - 64'd746842370399115, - 64'd240179086059323, - 64'd4887595867794, - 64'd626355321810053, - 64'd241323769247672, - 64'd9924776034165, - 64'd506183644970437, - 64'd239045080261808, - 64'd14449277222949, - 64'd387966088324595, - 64'd233629665829313, - 64'd18436722602651, - 64'd273192242411343, - 64'd225386198447957, - 64'd21871980748900, - 64'd163193051399847, - 64'd214639465259820, - 64'd24748685931934, - 64'd59134226199680, - 64'd201724674550048, - 64'd27068672904946, 64'd37987565983178, - 64'd186982042405970, - 64'd28841340383285, 64'd127345889852109, - 64'd170751713536614, - 64'd30082957333395, 64'd208283286974387, - 64'd153369061606049, - 64'd30815925929228, 64'd280307776928200, - 64'd135160405804480, - 64'd31068014600502, 64'd343087330259404, - 64'd116439171886633, - 64'd30871574010424, 64'd396442540850866, - 64'd97502517655162, - 64'd30262748079906, 64'd440337733251421, - 64'd78628434953589, - 64'd29280691340780, 64'd474870744605419, - 64'd60073332742995, - 64'd27966802972162, 64'd500261621297886, - 64'd42070098841254, - 64'd26363986871690, 64'd516840467547726, - 64'd24826631463055, - 64'd24515946056310, 64'd525034677232123, - 64'd8524825860936, - 64'd22466518594256, 64'd525355771520235, 64'd6680003832020, - 64'd20259061158714, 64'd518386053759184, 64'd20659291994046, - 64'd17935885181011, 64'd504765279825352, 64'd33311006438020, - 64'd15537749482665}};
	localparam logic signed[63:0] Fbi[0:2][0:74] = '{
		'{64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0, 64'd0},
		'{- 64'd459614617670948, 64'd236180802864224, 64'd53067997093561, - 64'd569532879783993, 64'd204301835870795, 64'd52855387393211, - 64'd663381517092044, 64'd171972686754111, 64'd51927510495402, - 64'd741059977026027, 64'd139674092112747, 64'd50350506447889, - 64'd802698871570680, 64'd107850538956602, 64'd48194565130026, - 64'd848640943034727, 64'd76906817930726, 64'd45532653550627, - 64'd879420514097390, 64'd47205382502847, 64'd42439299579991, - 64'd895741819343958, 64'd19064490578595, 64'd38989444734119, - 64'd898456601372454, - 64'd7242904060338, 64'd35257376733643, - 64'd888541336176843, - 64'd31489551041779, 64'd31315750657421, - 64'd867074430460488, - 64'd53493640748254, 64'd27234705627979, - 64'd835213708385532, - 64'd73117932686057, 64'd23081082127544, - 64'd794174477598151, - 64'd90268332318900, 64'd18917743271502, - 64'd745208434756558, - 64'd104891977155066, 64'd14803001680187, - 64'd689583639782946, - 64'd116974895134814, 64'd10790152006959, - 64'd628565756194885, - 64'd126539299582327, 64'd6927107714744, - 64'd563400722650966, - 64'd133640585224329, 64'd3256139356123, - 64'd495298988741795, - 64'd138364089105400, - 64'd186289587403, - 64'd425421416506145, - 64'd140821678725097, - 64'd3369594306864, - 64'd354866918548485, - 64'd141148227467154, - 64'd6269053615551, - 64'd284661874330815, - 64'd139498034473248, - 64'd8865714912952, - 64'd215751338517271, - 64'd136041242623042, - 64'd11146226438403, - 64'd148992029427446, - 64'd130960304309206, - 64'd13102604553515, - 64'd85147061921491, - 64'd124446540332005, - 64'd14731944114389, - 64'd24882367569355, - 64'd116696832572115, - 64'd16036080181081},
		'{64'd459614617670948, - 64'd236180802864224, - 64'd53067997093561, 64'd569532879783993, - 64'd204301835870795, - 64'd52855387393211, 64'd663381517092044, - 64'd171972686754111, - 64'd51927510495402, 64'd741059977026027, - 64'd139674092112747, - 64'd50350506447889, 64'd802698871570680, - 64'd107850538956602, - 64'd48194565130026, 64'd848640943034728, - 64'd76906817930726, - 64'd45532653550627, 64'd879420514097390, - 64'd47205382502847, - 64'd42439299579991, 64'd895741819343958, - 64'd19064490578595, - 64'd38989444734119, 64'd898456601372454, 64'd7242904060338, - 64'd35257376733643, 64'd888541336176843, 64'd31489551041779, - 64'd31315750657421, 64'd867074430460488, 64'd53493640748254, - 64'd27234705627979, 64'd835213708385532, 64'd73117932686057, - 64'd23081082127544, 64'd794174477598151, 64'd90268332318900, - 64'd18917743271502, 64'd745208434756558, 64'd104891977155066, - 64'd14803001680187, 64'd689583639782946, 64'd116974895134814, - 64'd10790152006959, 64'd628565756194885, 64'd126539299582327, - 64'd6927107714744, 64'd563400722650966, 64'd133640585224329, - 64'd3256139356123, 64'd495298988741795, 64'd138364089105400, 64'd186289587403, 64'd425421416506145, 64'd140821678725097, 64'd3369594306864, 64'd354866918548485, 64'd141148227467154, 64'd6269053615551, 64'd284661874330815, 64'd139498034473249, 64'd8865714912952, 64'd215751338517271, 64'd136041242623042, 64'd11146226438403, 64'd148992029427446, 64'd130960304309206, 64'd13102604553515, 64'd85147061921491, 64'd124446540332005, 64'd14731944114389, 64'd24882367569355, 64'd116696832572115, 64'd16036080181081}};
	localparam logic signed[63:0] hf[0:899] = {64'd11945802465280, - 64'd88788992000, - 64'd135408893952, 64'd11854973763584, - 64'd263853948928, - 64'd130432483328, 64'd11678164975616, - 64'd432925212672, - 64'd121096372224, 64'd11419062894592, - 64'd593334566912, - 64'd108066889728, 64'd11082592681984, - 64'd742788562944, - 64'd91996372992, 64'd10674729123840, - 64'd879368732672, - 64'd73516335104, 64'd10202312081408, - 64'd1001525805056, - 64'd53231304704, 64'd9672866136064, - 64'd1108070629376, - 64'd31713456128, 64'd9094416039936, - 64'd1198160084992, - 64'd9497970688, 64'd8475329429504, - 64'd1271280304128, 64'd12920766464, 64'd7824145907712, - 64'd1327226290176, 64'd35092201472, 64'd7149437059072, - 64'd1366078914560, 64'd56611872768, 64'd6459664891904, - 64'd1388180668416, 64'd77122895872, 64'd5763060203520, - 64'd1394108268544, 64'd96316768256, 64'd5067510382592, - 64'd1384646180864, 64'd113933434880, 64'd4380465299456, - 64'd1360757784576, 64'd129760763904, 64'd3708852895744, - 64'd1323556929536, 64'd143633432576, 64'd3059012861952, - 64'd1274279624704, 64'd155431256064, 64'd2436641062912, - 64'd1214256644096, 64'd165077057536, 64'd1846750740480, - 64'd1144886525952, 64'd172534169600, 64'd1293644333056, - 64'd1067609292800, 64'd177803542528, 64'd780898926592, - 64'd983883251712, 64'd180920598528, 64'd311363469312, - 64'd895161335808, 64'd181951873024, - 64'd112833470464, - 64'd802870984704, 64'd180991459328, - 64'd490266034176, - 64'd708394942464, 64'd178157404160, - 64'd820184285184, - 64'd613054808064, 64'd173588054016, - 64'd1102480015360, - 64'd518096453632, 64'd167438368768, - 64'd1337645465600, - 64'd424677507072, 64'd159876349952, - 64'd1526726524928, - 64'd333857226752, 64'd151079550976, - 64'd1671271677952, - 64'd246588620800, 64'd141231702016, - 64'd1773277020160, - 64'd163712516096, 64'd130519572480, - 64'd1835129372672, - 64'd85953642496, 64'd119129956352, - 64'd1859547299840, - 64'd13918779392, 64'd107246985216, - 64'd1849522782208, 64'd51903332352, 64'd95049629696, - 64'd1808261709824, 64'd111140438016, 64'd82709463040, - 64'd1739127128064, 64'd163533651968, 64'd70388752384, - 64'd1645583007744, 64'd208932978688, 64'd58238791680, - 64'd1531141947392, 64'd247291691008, 64'd46398500864, - 64'd1399314448384, 64'd278659530752, 64'd34993369088, - 64'd1253563301888, 64'd303175204864, 64'd24134610944, - 64'd1097260859392, 64'd321058177024, 64'd13918623744, - 64'd933651021824, 64'd332599754752, 64'd4426675712, - 64'd765815422976, 64'd338154061824, - 64'd4275155712, - 64'd596644790272, 64'd338128666624, - 64'd12135829504, - 64'd428814368768, 64'd332975144960, - 64'd19118987264, - 64'd264764375040, 64'd323179839488, - 64'd25202413568, - 64'd106685071360, 64'd309254619136, - 64'd30377345024, 64'd43493859328, 64'd291728162816, - 64'd34647633920, 64'd184109432832, 64'd271137488896, - 64'd38028791808, 64'd313767526400, 64'd248020058112, - 64'd40546959360, 64'd431341273088, 64'd222906515456, - 64'd42237788160, 64'd535965761536, 64'd196313890816, - 64'd43145261056, 64'd627029770240, 64'd168739651584, - 64'd43320508416, 64'd704164528128, 64'd140656345088, - 64'd42820591616, 64'd767230214144, 64'd112507068416, - 64'd41707307008, 64'd816299966464, 64'd84701552640, - 64'd40045989888, 64'd851642548224, 64'd57613160448, - 64'd37904388096, 64'd873703669760, 64'd31576444928, - 64'd35351556096, 64'd883085672448, 64'd6885519872, - 64'd32456830976, 64'd880527605760, - 64'd16206928896, - 64'd29288859648, 64'd866883993600, - 64'd37489987584, - 64'd25914730496, 64'd843104124928, - 64'd56794263552, - 64'd22399170560, 64'd810211672064, - 64'd73991069696, - 64'd18803847168, 64'd769284243456, - 64'd88991121408, - 64'd15186750464, 64'd721434509312, - 64'd101742788608, - 64'd11601685504, 64'd667791785984, - 64'd112229965824, - 64'd8097846784, 64'd609484734464, - 64'd120469594112, - 64'd4719493632, 64'd547625828352, - 64'd126508924928, - 64'd1505719424, 64'd483296739328, - 64'd130422595584, 64'd1509698176, 64'd417535459328, - 64'd132309491712, 64'd4298357248, 64'd351325093888, - 64'd132289552384, 64'd6837216768, 64'd285584097280, - 64'd130500534272, 64'd9108505600, 64'd221158211584, - 64'd127094710272, 64'd11099573248, 64'd158814011392, - 64'd122235699200, 64'd12802669568, 64'd99234119680, - 64'd116095311872, 64'd14214686720, 64'd43013812224, - 64'd108850552832, 64'd15336848384, - 64'd9340810240, - 64'd100680744960, 64'd16174363648, - 64'd57413300224, - 64'd91764891648, 64'd16736053248, - 64'd100876050432, - 64'd82279178240, 64'd17033956352, - 64'd139488313344, - 64'd72394743808, 64'd17082915840, - 64'd173093142528, - 64'd62275670016, 64'd16900162560, - 64'd201613426688, - 64'd52077232128, 64'd16504897536, - 64'd225047052288, - 64'd41944383488, 64'd15917870080, - 64'd243461505024, - 64'd32010526720, 64'd15160978432, - 64'd256987693056, - 64'd22396487680, 64'd14256874496, - 64'd265813573632, - 64'd13209807872, 64'd13228594176, - 64'd270177353728, - 64'd4544207360, 64'd12099204096, - 64'd270360428544, 64'd3520669952, 64'd10891482112, - 64'd266680434688, 64'd10919326720, 64'd9627619328, - 64'd259484123136, 64'd17600268288, 64'd8328953856, - 64'd249140477952, 64'd23525679104, 64'd7015740416, - 64'd236033982464, 64'd28670932992, 64'd5706946560, - 64'd220558147584, 64'd33023950848, 64'd4420085760, - 64'd203109548032, 64'd36584452096, 64'd3171081728, - 64'd184081989632, 64'd39363063808, 64'd1974165376, - 64'd163861413888, 64'd41380384768, 64'd841802944, - 64'd142821130240, 64'd42665955328, - 64'd215346240, - 64'd121317605376, 64'd43257176064, - 64'd1188443648, - 64'd99686866944, 64'd43198226432, - 64'd2070459264, - 64'd78241341440, 64'd42538938368, - 64'd2856134400, - 64'd57267331072, 64'd41333694464, - 64'd3541924096, - 64'd37023051776, 64'd39640338432, - 64'd4125918464, - 64'd17737127936, 64'd37519114240, - 64'd4607749120, 64'd392314560, 64'd35031670784, - 64'd4988478464, 64'd17198120960, 64'd32240097280, - 64'd5270480896, 64'd32544086016, 64'd29206026240, - 64'd5457310720, 64'd46324523008, 64'd25989832704, - 64'd5553567744, 64'd58463432704, 64'd22649884672, - 64'd5564754944, 64'd68913340416, 64'd19241889792, - 64'd5497134592, 64'd77653811200, 64'd15818323968, - 64'd5357588992, 64'd84689698816, 64'd12427952128, - 64'd5153475072, 64'd90049191936, 64'd9115423744, - 64'd4892490240, 64'd93781688320, 64'd5920968192, - 64'd4582541824, 64'd95955509248, 64'd2880170496, - 64'd4231618816, 64'd96655523840, 64'd23821962, - 64'd3847678976, 64'd95980765184, - 64'd2622145024, - 64'd3438540032, 64'd94041980928, - 64'd5036652544, - 64'd3011781888, 64'd90959224832, - 64'd7203406336, - 64'd2574660096, 64'd86859497472, - 64'd9110765568, - 64'd2134030848, 64'd81874468864, - 64'd10751552512, - 64'd1696284160, 64'd76138291200, - 64'd12122821632, - 64'd1267292160, 64'd69785583616, - 64'd13225584640, - 64'd852365568, 64'd62949490688, - 64'd14064497664, - 64'd456222880, 64'd55759986688, - 64'd14647527424, - 64'd82969016, 64'd48342290432, - 64'd14985594880, 64'd263915376, 64'd40815476736, - 64'd15092198400, 64'd581575552, 64'd33291302912, - 64'd14983040000, 64'd867775296, 64'd25873192960, - 64'd14675641344, 64'd1120881792, 64'd18655430656, - 64'd14188963840, 64'd1339842816, 64'd11722529792, - 64'd13543043072, 64'd1524158208, 64'd5148798464, - 64'd12758625280, 64'd1673845632, - 64'd1001938752, - 64'd11856831488, 64'd1789401344, - 64'd6676438528, - 64'd10858838016, 64'd1871757824, - 64'd11831991296, - 64'd9785572352, 64'd1922238080, - 64'd16436226048, - 64'd8657452032, 64'd1942508416, - 64'd20466792448, - 64'd7494131200, 64'd1934529664, - 64'd23910922240, - 64'd6314289664, 64'd1900507904, - 64'd26764894208, - 64'd5135446528, 64'd1842845824, - 64'd29033412608, - 64'd3973803776, 64'd1764094592, - 64'd30728910848, - 64'd2844120064, 64'd1666907776, - 64'd31870814208, - 64'd1759613696, 64'd1553996416, - 64'd32484743168, - 64'd731895616, 64'd1428087680, - 64'd32601698304, 64'd229072928, 64'd1291885824, - 64'd32257234944, 64'd1114994432, 64'd1148036352, - 64'd31490633728, 64'd1919226496, 64'd999093824, - 64'd30344075264, 64'd2636750336, 64'd847493056, - 64'd28861843456, 64'd3264119040, 64'd695524800, - 64'd27089559552, 64'd3799388928, 64'd545314240, - 64'd25073446912, 64'd4242033408, 64'd398804416, - 64'd22859651072, 64'd4592845824, 64'd257742464, - 64'd20493606912, 64'd4853829632, 64'd123670304, - 64'd18019463168, 64'd5028080640, - 64'd2081519, - 64'd15479568384, 64'd5119662080, - 64'd118396488, - 64'd12914020352, 64'd5133478400, - 64'd224371632, - 64'd10360278016, 64'd5075143168, - 64'd319314080, - 64'd7852839424, 64'd4950847488, - 64'd402735040, - 64'd5422990336, 64'd4767235584, - 64'd474341376, - 64'd3098605312, 64'd4531273728, - 64'd534025024, - 64'd904020672, 64'd4250134272, - 64'd581850816, 64'd1140039808, 64'd3931079168, - 64'd618042496, 64'd3016482048, 64'd3581352704, - 64'd642968128, 64'd4711806976, 64'd3208083968, - 64'd657124032, 64'd6216029696, 64'd2818194944, - 64'd661118208, 64'd7522554880, 64'd2418322432, - 64'd655654080, 64'd8628016128, 64'd2014745472, - 64'd641513152, 64'd9532080128, 64'd1613326592, - 64'd619538880, 64'd10237225984, 64'd1219460992, - 64'd590619840, 64'd10748503040, 64'd838037376, - 64'd555674624, 64'd11073265664, 64'd473407520, - 64'd515636544, 64'd11220903936, 64'd129366392, - 64'd471439744, 64'd11202555904, - 64'd190858784, - 64'd424006240, 64'd11030830080, - 64'd484610944, - 64'd374234016, 64'd10719516672, - 64'd749797440, - 64'd322986496, 64'd10283310080, - 64'd984876800, - 64'd271083072, 64'd9737539584, - 64'd1188839168, - 64'd219291104, 64'd9097907200, - 64'd1361180288, - 64'd168319184, 64'd8380242944, - 64'd1501871360, - 64'd118811752, 64'd7600279552, - 64'd1611323264, - 64'd71344880, 64'd6773438976, - 64'd1690348672, - 64'd26423486, 64'd5914642432, - 64'd1740120832, 64'd15520401, 64'd5038141952, - 64'd1762129920, 64'd54128152, 64'd4157373696, - 64'd1758139392, 64'd89114032, 64'd3284831232, - 64'd1730141056, 64'd120263744, 64'd2431964160, - 64'd1680310400, 64'd147432016, 64'd1609096832, - 64'd1610962816, 64'd170539504, 64'd825370176, - 64'd1524511104, 64'd189568992, 64'd88702496, - 64'd1423424896, 64'd204560944, - 64'd594228416, - 64'd1310192512, 64'd215608672, - 64'd1217985280, - 64'd1187284608, 64'd222853120, - 64'd1778354560, - 64'd1057121792, 64'd226477344, - 64'd2272312832, - 64'd922044544, 64'd226700864, - 64'd2697980416, - 64'd784286976, 64'd223773840, - 64'd3054562304, - 64'd645953920, 64'd217971456, - 64'd3342277632, - 64'd509001120, 64'd209588096, - 64'd3562282240, - 64'd375219744, 64'd198931952, - 64'd3716581632, - 64'd246223504, 64'd186319712, - 64'd3807940608, - 64'd123439736, 64'd172071488, - 64'd3839788544, - 64'd8103470, 64'd156506192, - 64'd3816122112, 64'd98745264, 64'd139937200, - 64'd3741408000, 64'd196261344, 64'd122668424, - 64'd3620485888, 64'd283791712, 64'd104990800, - 64'd3458473472, 64'd360870016, 64'd87179240, - 64'd3260676096, 64'd427209344, 64'd69490048, - 64'd3032497664, 64'd482692544, 64'd52158712, - 64'd2779360256, 64'd527361472, 64'd35398248, - 64'd2506626816, 64'd561404352, 64'd19397894, - 64'd2219531008, 64'd585142336, 64'd4322274, - 64'd1923115776, 64'd599015296, - 64'd9689042, - 64'd1622176640, 64'd603566656, - 64'd22521606, - 64'd1321214592, 64'd599428288, - 64'd34085796, - 64'd1024395072, 64'd587305152, - 64'd44316220, - 64'd735515904, 64'd567960128, - 64'd53170792, - 64'd457981920, 64'd542199168, - 64'd60629608, - 64'd194787280, 64'd510856832, - 64'd66693536, 64'd51495420, 64'd474782720, - 64'd71382688, 64'd278719296, 64'd434828512, - 64'd74734672, 64'd485161088, 64'd391836160, - 64'd76802800, 64'd669513536, 64'd346626816, - 64'd77654168, 64'd830872320, 64'd299991136, - 64'd77367704, 64'd968718656, 64'd252680544, - 64'd76032176, 64'd1082897664, 64'd205399824, - 64'd73744264, 64'd1173593344, 64'd158800832, - 64'd70606600, 64'd1241300992, 64'd113477360, - 64'd66725936, 64'd1286796928, 64'd69961344, - 64'd62211332, 64'd1311106816, 64'd28720044, - 64'd57172488, 64'd1315473024, - 64'd9845552, - 64'd51718192, 64'd1301321088, - 64'd45401364, - 64'd45954856, 64'd1270226688, - 64'd77679840, - 64'd39985240, 64'd1223882368, - 64'd106478696, - 64'd33907308, 64'd1164065536, - 64'd131658880, - 64'd27813206, 64'd1092607232, - 64'd153141728, - 64'd21788444, 64'd1011363392, - 64'd170905616, - 64'd15911199, 64'd922186944, - 64'd184981952, - 64'd10251780, 64'd826902336, - 64'd195450800, - 64'd4872242, 64'd727282752, - 64'd202436224, 64'd173855, 64'd625029056, - 64'd206101136, 64'd4841557, 64'd521751808, - 64'd206642320, 64'd9094493, 64'd418955744, - 64'd204285040, 64'd12904741, 64'd318026816, - 64'd199277920, 64'd16252584, 64'd220221824, - 64'd191887664, 64'd19126170, 64'd126660776, - 64'd182394096, 64'd21521090, 64'd38321452, - 64'd171085264, 64'd23439886, - 64'd43963440, - 64'd158252880, 64'd24891498, - 64'd119506984, - 64'd144187968, 64'd25890662, - 64'd187766720, - 64'd129176920, 64'd26457268, - 64'd248341328, - 64'd113497880, 64'd26615718, - 64'd300965728, - 64'd97417504, 64'd26394232, - 64'd345504544, - 64'd81188104, 64'd25824188, - 64'd381944352, - 64'd65045288, 64'd24939446, - 64'd410384704, - 64'd49205876, 64'd23775694, - 64'd431028384, - 64'd33866352, 64'd22369818, - 64'd444171008, - 64'd19201632, 64'd20759312, - 64'd450189760, - 64'd5364273, 64'd18981700, - 64'd449532352, 64'd7515990, 64'd17074022, - 64'd442705472, 64'd19332324, 64'd15072356, - 64'd430263360, 64'd30000578, 64'd13011396, - 64'd412796608, 64'd39458748, 64'd10924065, - 64'd390921312, 64'd47666192, 64'd8841202, - 64'd365268608, 64'd54602596, 64'd6791282, - 64'd336474912, 64'd60266744, 64'd4800206, - 64'd305172576, 64'd64675104, 64'd2891127, - 64'd271981568, 64'd67860288, 64'd1084341, - 64'd237501760, 64'd69869392, - 64'd602783, - 64'd202306160, 64'd70762288, - 64'd2155828, - 64'd166934976, 64'd70609800, - 64'd3563304, - 64'd131890544, 64'd69491960, - 64'd4816591, - 64'd97633288, 64'd67496168, - 64'd5909846, - 64'd64578416, 64'd64715456, - 64'd6839872, - 64'd33093550, 64'd61246792, - 64'd7605972, - 64'd3497204, 64'd57189428, - 64'd8209764, 64'd23941968, 64'd52643360, - 64'd8654994, 64'd49005176, 64'd47707892, - 64'd8947319, 64'd71522792, 64'd42480312, - 64'd9094092, 64'd91373056, 64'd37054708, - 64'd9104131, 64'd108480168, 64'd31520876, - 64'd8987487, 64'd122811920, 64'd25963438, - 64'd8755215, 64'd134376896, 64'd20461020, - 64'd8419144, 64'd143221328, 64'd15085639, - 64'd7991660, 64'd149425616, 64'd9902178, - 64'd7485490, 64'd153100688, 64'd4968036, - 64'd6913496, 64'd154384208, 64'd332884, - 64'd6288499, 64'd153436624, - 64'd3961446, - 64'd5623094, 64'd150437328, - 64'd7880952, - 64'd4929494, 64'd145580704, - 64'd11399351, - 64'd4219398, 64'd139072352, - 64'd14497869, - 64'd3503856, 64'd131125376, - 64'd17164936, - 64'd2793172, 64'd121956920, - 64'd19395814, - 64'd2096814, 64'd111784840, - 64'd21192152, - 64'd1423346, 64'd100824616, - 64'd22561486, - 64'd780380, 64'd89286600, - 64'd23516698, - 64'd174535, 64'd77373448, - 64'd24075436, 64'd388574, 64'd65277892, - 64'd24259520, 64'd904344, 64'd53180840, - 64'd24094322, 64'd1369168, 64'd41249728, - 64'd23608160, 64'd1780413, 64'd29637228, - 64'd22831676, 64'd2136383, 64'd18480216, - 64'd21797248, 64'd2436275, 64'd7899076, - 64'd20538406, 64'd2680118, - 64'd2002750, - 64'd19089290, 64'd2868718, - 64'd11138924, - 64'd17484122, 64'd3003581, - 64'd19440132, - 64'd15756735, 64'd3086848};
	localparam logic signed[63:0] hb[0:899] = {64'd11945802465280, 64'd88788992000, - 64'd135408893952, 64'd11854973763584, 64'd263853948928, - 64'd130432483328, 64'd11678164975616, 64'd432925212672, - 64'd121096372224, 64'd11419062894592, 64'd593334566912, - 64'd108066889728, 64'd11082592681984, 64'd742788562944, - 64'd91996372992, 64'd10674729123840, 64'd879368732672, - 64'd73516335104, 64'd10202312081408, 64'd1001525805056, - 64'd53231304704, 64'd9672866136064, 64'd1108070629376, - 64'd31713456128, 64'd9094416039936, 64'd1198160084992, - 64'd9497970688, 64'd8475329429504, 64'd1271280304128, 64'd12920766464, 64'd7824145907712, 64'd1327226290176, 64'd35092201472, 64'd7149437059072, 64'd1366078914560, 64'd56611872768, 64'd6459664891904, 64'd1388180668416, 64'd77122895872, 64'd5763060203520, 64'd1394108268544, 64'd96316768256, 64'd5067510382592, 64'd1384646180864, 64'd113933434880, 64'd4380465299456, 64'd1360757784576, 64'd129760763904, 64'd3708852895744, 64'd1323556929536, 64'd143633432576, 64'd3059012861952, 64'd1274279624704, 64'd155431256064, 64'd2436641062912, 64'd1214256644096, 64'd165077057536, 64'd1846750740480, 64'd1144886525952, 64'd172534169600, 64'd1293644333056, 64'd1067609292800, 64'd177803542528, 64'd780898926592, 64'd983883251712, 64'd180920598528, 64'd311363469312, 64'd895161335808, 64'd181951873024, - 64'd112833470464, 64'd802870984704, 64'd180991459328, - 64'd490266034176, 64'd708394942464, 64'd178157404160, - 64'd820184285184, 64'd613054808064, 64'd173588054016, - 64'd1102480015360, 64'd518096453632, 64'd167438368768, - 64'd1337645465600, 64'd424677507072, 64'd159876349952, - 64'd1526726524928, 64'd333857226752, 64'd151079550976, - 64'd1671271677952, 64'd246588620800, 64'd141231702016, - 64'd1773277020160, 64'd163712516096, 64'd130519572480, - 64'd1835129372672, 64'd85953642496, 64'd119129956352, - 64'd1859547299840, 64'd13918779392, 64'd107246985216, - 64'd1849522782208, - 64'd51903332352, 64'd95049629696, - 64'd1808261709824, - 64'd111140438016, 64'd82709463040, - 64'd1739127128064, - 64'd163533651968, 64'd70388752384, - 64'd1645583007744, - 64'd208932978688, 64'd58238791680, - 64'd1531141947392, - 64'd247291691008, 64'd46398500864, - 64'd1399314448384, - 64'd278659530752, 64'd34993369088, - 64'd1253563301888, - 64'd303175204864, 64'd24134610944, - 64'd1097260859392, - 64'd321058177024, 64'd13918623744, - 64'd933651021824, - 64'd332599754752, 64'd4426675712, - 64'd765815422976, - 64'd338154061824, - 64'd4275155712, - 64'd596644790272, - 64'd338128666624, - 64'd12135829504, - 64'd428814368768, - 64'd332975144960, - 64'd19118987264, - 64'd264764375040, - 64'd323179839488, - 64'd25202413568, - 64'd106685071360, - 64'd309254619136, - 64'd30377345024, 64'd43493859328, - 64'd291728162816, - 64'd34647633920, 64'd184109432832, - 64'd271137488896, - 64'd38028791808, 64'd313767526400, - 64'd248020058112, - 64'd40546959360, 64'd431341273088, - 64'd222906515456, - 64'd42237788160, 64'd535965761536, - 64'd196313890816, - 64'd43145261056, 64'd627029770240, - 64'd168739651584, - 64'd43320508416, 64'd704164528128, - 64'd140656345088, - 64'd42820591616, 64'd767230214144, - 64'd112507068416, - 64'd41707307008, 64'd816299966464, - 64'd84701552640, - 64'd40045989888, 64'd851642548224, - 64'd57613160448, - 64'd37904388096, 64'd873703669760, - 64'd31576444928, - 64'd35351556096, 64'd883085672448, - 64'd6885519872, - 64'd32456830976, 64'd880527605760, 64'd16206928896, - 64'd29288859648, 64'd866883993600, 64'd37489987584, - 64'd25914730496, 64'd843104124928, 64'd56794263552, - 64'd22399170560, 64'd810211672064, 64'd73991069696, - 64'd18803847168, 64'd769284243456, 64'd88991121408, - 64'd15186750464, 64'd721434509312, 64'd101742788608, - 64'd11601685504, 64'd667791785984, 64'd112229965824, - 64'd8097846784, 64'd609484734464, 64'd120469594112, - 64'd4719493632, 64'd547625828352, 64'd126508924928, - 64'd1505719424, 64'd483296739328, 64'd130422595584, 64'd1509698176, 64'd417535459328, 64'd132309491712, 64'd4298357248, 64'd351325093888, 64'd132289552384, 64'd6837216768, 64'd285584097280, 64'd130500534272, 64'd9108505600, 64'd221158211584, 64'd127094710272, 64'd11099573248, 64'd158814011392, 64'd122235699200, 64'd12802669568, 64'd99234119680, 64'd116095311872, 64'd14214686720, 64'd43013812224, 64'd108850552832, 64'd15336848384, - 64'd9340810240, 64'd100680744960, 64'd16174363648, - 64'd57413300224, 64'd91764891648, 64'd16736053248, - 64'd100876050432, 64'd82279178240, 64'd17033956352, - 64'd139488313344, 64'd72394743808, 64'd17082915840, - 64'd173093142528, 64'd62275670016, 64'd16900162560, - 64'd201613426688, 64'd52077232128, 64'd16504897536, - 64'd225047052288, 64'd41944383488, 64'd15917870080, - 64'd243461505024, 64'd32010526720, 64'd15160978432, - 64'd256987693056, 64'd22396487680, 64'd14256874496, - 64'd265813573632, 64'd13209807872, 64'd13228594176, - 64'd270177353728, 64'd4544207360, 64'd12099204096, - 64'd270360428544, - 64'd3520669952, 64'd10891482112, - 64'd266680434688, - 64'd10919326720, 64'd9627619328, - 64'd259484123136, - 64'd17600268288, 64'd8328953856, - 64'd249140477952, - 64'd23525679104, 64'd7015740416, - 64'd236033982464, - 64'd28670932992, 64'd5706946560, - 64'd220558147584, - 64'd33023950848, 64'd4420085760, - 64'd203109548032, - 64'd36584452096, 64'd3171081728, - 64'd184081989632, - 64'd39363063808, 64'd1974165376, - 64'd163861413888, - 64'd41380384768, 64'd841802944, - 64'd142821130240, - 64'd42665955328, - 64'd215346240, - 64'd121317605376, - 64'd43257176064, - 64'd1188443648, - 64'd99686866944, - 64'd43198226432, - 64'd2070459264, - 64'd78241341440, - 64'd42538938368, - 64'd2856134400, - 64'd57267331072, - 64'd41333694464, - 64'd3541924096, - 64'd37023051776, - 64'd39640338432, - 64'd4125918464, - 64'd17737127936, - 64'd37519114240, - 64'd4607749120, 64'd392314560, - 64'd35031670784, - 64'd4988478464, 64'd17198120960, - 64'd32240097280, - 64'd5270480896, 64'd32544086016, - 64'd29206026240, - 64'd5457310720, 64'd46324523008, - 64'd25989832704, - 64'd5553567744, 64'd58463432704, - 64'd22649884672, - 64'd5564754944, 64'd68913340416, - 64'd19241889792, - 64'd5497134592, 64'd77653811200, - 64'd15818323968, - 64'd5357588992, 64'd84689698816, - 64'd12427952128, - 64'd5153475072, 64'd90049191936, - 64'd9115423744, - 64'd4892490240, 64'd93781688320, - 64'd5920968192, - 64'd4582541824, 64'd95955509248, - 64'd2880170496, - 64'd4231618816, 64'd96655523840, - 64'd23821962, - 64'd3847678976, 64'd95980765184, 64'd2622145024, - 64'd3438540032, 64'd94041980928, 64'd5036652544, - 64'd3011781888, 64'd90959224832, 64'd7203406336, - 64'd2574660096, 64'd86859497472, 64'd9110765568, - 64'd2134030848, 64'd81874468864, 64'd10751552512, - 64'd1696284160, 64'd76138291200, 64'd12122821632, - 64'd1267292160, 64'd69785583616, 64'd13225584640, - 64'd852365568, 64'd62949490688, 64'd14064497664, - 64'd456222880, 64'd55759986688, 64'd14647527424, - 64'd82969016, 64'd48342290432, 64'd14985594880, 64'd263915376, 64'd40815476736, 64'd15092198400, 64'd581575552, 64'd33291302912, 64'd14983040000, 64'd867775296, 64'd25873192960, 64'd14675641344, 64'd1120881792, 64'd18655430656, 64'd14188963840, 64'd1339842816, 64'd11722529792, 64'd13543043072, 64'd1524158208, 64'd5148798464, 64'd12758625280, 64'd1673845632, - 64'd1001938752, 64'd11856831488, 64'd1789401344, - 64'd6676438528, 64'd10858838016, 64'd1871757824, - 64'd11831991296, 64'd9785572352, 64'd1922238080, - 64'd16436226048, 64'd8657452032, 64'd1942508416, - 64'd20466792448, 64'd7494131200, 64'd1934529664, - 64'd23910922240, 64'd6314289664, 64'd1900507904, - 64'd26764894208, 64'd5135446528, 64'd1842845824, - 64'd29033412608, 64'd3973803776, 64'd1764094592, - 64'd30728910848, 64'd2844120064, 64'd1666907776, - 64'd31870814208, 64'd1759613696, 64'd1553996416, - 64'd32484743168, 64'd731895616, 64'd1428087680, - 64'd32601698304, - 64'd229072928, 64'd1291885824, - 64'd32257234944, - 64'd1114994432, 64'd1148036352, - 64'd31490633728, - 64'd1919226496, 64'd999093824, - 64'd30344075264, - 64'd2636750336, 64'd847493056, - 64'd28861843456, - 64'd3264119040, 64'd695524800, - 64'd27089559552, - 64'd3799388928, 64'd545314240, - 64'd25073446912, - 64'd4242033408, 64'd398804416, - 64'd22859651072, - 64'd4592845824, 64'd257742464, - 64'd20493606912, - 64'd4853829632, 64'd123670304, - 64'd18019463168, - 64'd5028080640, - 64'd2081519, - 64'd15479568384, - 64'd5119662080, - 64'd118396488, - 64'd12914020352, - 64'd5133478400, - 64'd224371632, - 64'd10360278016, - 64'd5075143168, - 64'd319314080, - 64'd7852839424, - 64'd4950847488, - 64'd402735040, - 64'd5422990336, - 64'd4767235584, - 64'd474341376, - 64'd3098605312, - 64'd4531273728, - 64'd534025024, - 64'd904020672, - 64'd4250134272, - 64'd581850816, 64'd1140039808, - 64'd3931079168, - 64'd618042496, 64'd3016482048, - 64'd3581352704, - 64'd642968128, 64'd4711806976, - 64'd3208083968, - 64'd657124032, 64'd6216029696, - 64'd2818194944, - 64'd661118208, 64'd7522554880, - 64'd2418322432, - 64'd655654080, 64'd8628016128, - 64'd2014745472, - 64'd641513152, 64'd9532080128, - 64'd1613326592, - 64'd619538880, 64'd10237225984, - 64'd1219460992, - 64'd590619840, 64'd10748503040, - 64'd838037376, - 64'd555674624, 64'd11073265664, - 64'd473407520, - 64'd515636544, 64'd11220903936, - 64'd129366392, - 64'd471439744, 64'd11202555904, 64'd190858784, - 64'd424006240, 64'd11030830080, 64'd484610944, - 64'd374234016, 64'd10719516672, 64'd749797440, - 64'd322986496, 64'd10283310080, 64'd984876800, - 64'd271083072, 64'd9737539584, 64'd1188839168, - 64'd219291104, 64'd9097907200, 64'd1361180288, - 64'd168319184, 64'd8380242944, 64'd1501871360, - 64'd118811752, 64'd7600279552, 64'd1611323264, - 64'd71344880, 64'd6773438976, 64'd1690348672, - 64'd26423486, 64'd5914642432, 64'd1740120832, 64'd15520401, 64'd5038141952, 64'd1762129920, 64'd54128152, 64'd4157373696, 64'd1758139392, 64'd89114032, 64'd3284831232, 64'd1730141056, 64'd120263744, 64'd2431964160, 64'd1680310400, 64'd147432016, 64'd1609096832, 64'd1610962816, 64'd170539504, 64'd825370176, 64'd1524511104, 64'd189568992, 64'd88702496, 64'd1423424896, 64'd204560944, - 64'd594228416, 64'd1310192512, 64'd215608672, - 64'd1217985280, 64'd1187284608, 64'd222853120, - 64'd1778354560, 64'd1057121792, 64'd226477344, - 64'd2272312832, 64'd922044544, 64'd226700864, - 64'd2697980416, 64'd784286976, 64'd223773840, - 64'd3054562304, 64'd645953920, 64'd217971456, - 64'd3342277632, 64'd509001120, 64'd209588096, - 64'd3562282240, 64'd375219744, 64'd198931952, - 64'd3716581632, 64'd246223504, 64'd186319712, - 64'd3807940608, 64'd123439736, 64'd172071488, - 64'd3839788544, 64'd8103470, 64'd156506192, - 64'd3816122112, - 64'd98745264, 64'd139937200, - 64'd3741408000, - 64'd196261344, 64'd122668424, - 64'd3620485888, - 64'd283791712, 64'd104990800, - 64'd3458473472, - 64'd360870016, 64'd87179240, - 64'd3260676096, - 64'd427209344, 64'd69490048, - 64'd3032497664, - 64'd482692544, 64'd52158712, - 64'd2779360256, - 64'd527361472, 64'd35398248, - 64'd2506626816, - 64'd561404352, 64'd19397894, - 64'd2219531008, - 64'd585142336, 64'd4322274, - 64'd1923115776, - 64'd599015296, - 64'd9689042, - 64'd1622176640, - 64'd603566656, - 64'd22521606, - 64'd1321214592, - 64'd599428288, - 64'd34085796, - 64'd1024395072, - 64'd587305152, - 64'd44316220, - 64'd735515904, - 64'd567960128, - 64'd53170792, - 64'd457981920, - 64'd542199168, - 64'd60629608, - 64'd194787280, - 64'd510856832, - 64'd66693536, 64'd51495420, - 64'd474782720, - 64'd71382688, 64'd278719296, - 64'd434828512, - 64'd74734672, 64'd485161088, - 64'd391836160, - 64'd76802800, 64'd669513536, - 64'd346626816, - 64'd77654168, 64'd830872320, - 64'd299991136, - 64'd77367704, 64'd968718656, - 64'd252680544, - 64'd76032176, 64'd1082897664, - 64'd205399824, - 64'd73744264, 64'd1173593344, - 64'd158800832, - 64'd70606600, 64'd1241300992, - 64'd113477360, - 64'd66725936, 64'd1286796928, - 64'd69961344, - 64'd62211332, 64'd1311106816, - 64'd28720044, - 64'd57172488, 64'd1315473024, 64'd9845552, - 64'd51718192, 64'd1301321088, 64'd45401364, - 64'd45954856, 64'd1270226688, 64'd77679840, - 64'd39985240, 64'd1223882368, 64'd106478696, - 64'd33907308, 64'd1164065536, 64'd131658880, - 64'd27813206, 64'd1092607232, 64'd153141728, - 64'd21788444, 64'd1011363392, 64'd170905616, - 64'd15911199, 64'd922186944, 64'd184981952, - 64'd10251780, 64'd826902336, 64'd195450800, - 64'd4872242, 64'd727282752, 64'd202436224, 64'd173855, 64'd625029056, 64'd206101136, 64'd4841557, 64'd521751808, 64'd206642320, 64'd9094493, 64'd418955744, 64'd204285040, 64'd12904741, 64'd318026816, 64'd199277920, 64'd16252584, 64'd220221824, 64'd191887664, 64'd19126170, 64'd126660776, 64'd182394096, 64'd21521090, 64'd38321452, 64'd171085264, 64'd23439886, - 64'd43963440, 64'd158252880, 64'd24891498, - 64'd119506984, 64'd144187968, 64'd25890662, - 64'd187766720, 64'd129176920, 64'd26457268, - 64'd248341328, 64'd113497880, 64'd26615718, - 64'd300965728, 64'd97417504, 64'd26394232, - 64'd345504544, 64'd81188104, 64'd25824188, - 64'd381944352, 64'd65045288, 64'd24939446, - 64'd410384704, 64'd49205876, 64'd23775694, - 64'd431028384, 64'd33866352, 64'd22369818, - 64'd444171008, 64'd19201632, 64'd20759312, - 64'd450189760, 64'd5364273, 64'd18981700, - 64'd449532352, - 64'd7515990, 64'd17074022, - 64'd442705472, - 64'd19332324, 64'd15072356, - 64'd430263360, - 64'd30000578, 64'd13011396, - 64'd412796608, - 64'd39458748, 64'd10924065, - 64'd390921312, - 64'd47666192, 64'd8841202, - 64'd365268608, - 64'd54602596, 64'd6791282, - 64'd336474912, - 64'd60266744, 64'd4800206, - 64'd305172576, - 64'd64675104, 64'd2891127, - 64'd271981568, - 64'd67860288, 64'd1084341, - 64'd237501760, - 64'd69869392, - 64'd602783, - 64'd202306160, - 64'd70762288, - 64'd2155828, - 64'd166934976, - 64'd70609800, - 64'd3563304, - 64'd131890544, - 64'd69491960, - 64'd4816591, - 64'd97633288, - 64'd67496168, - 64'd5909846, - 64'd64578416, - 64'd64715456, - 64'd6839872, - 64'd33093550, - 64'd61246792, - 64'd7605972, - 64'd3497204, - 64'd57189428, - 64'd8209764, 64'd23941968, - 64'd52643360, - 64'd8654994, 64'd49005176, - 64'd47707892, - 64'd8947319, 64'd71522792, - 64'd42480312, - 64'd9094092, 64'd91373056, - 64'd37054708, - 64'd9104131, 64'd108480168, - 64'd31520876, - 64'd8987487, 64'd122811920, - 64'd25963438, - 64'd8755215, 64'd134376896, - 64'd20461020, - 64'd8419144, 64'd143221328, - 64'd15085639, - 64'd7991660, 64'd149425616, - 64'd9902178, - 64'd7485490, 64'd153100688, - 64'd4968036, - 64'd6913496, 64'd154384208, - 64'd332884, - 64'd6288499, 64'd153436624, 64'd3961446, - 64'd5623094, 64'd150437328, 64'd7880952, - 64'd4929494, 64'd145580704, 64'd11399351, - 64'd4219398, 64'd139072352, 64'd14497869, - 64'd3503856, 64'd131125376, 64'd17164936, - 64'd2793172, 64'd121956920, 64'd19395814, - 64'd2096814, 64'd111784840, 64'd21192152, - 64'd1423346, 64'd100824616, 64'd22561486, - 64'd780380, 64'd89286600, 64'd23516698, - 64'd174535, 64'd77373448, 64'd24075436, 64'd388574, 64'd65277892, 64'd24259520, 64'd904344, 64'd53180840, 64'd24094322, 64'd1369168, 64'd41249728, 64'd23608160, 64'd1780413, 64'd29637228, 64'd22831676, 64'd2136383, 64'd18480216, 64'd21797248, 64'd2436275, 64'd7899076, 64'd20538406, 64'd2680118, - 64'd2002750, 64'd19089290, 64'd2868718, - 64'd11138924, 64'd17484122, 64'd3003581, - 64'd19440132, 64'd15756735, 64'd3086848};
endpackage
`endif
