`ifndef COEFFICIENTS_FX_SV_
`define COEFFICIENTS_FX_SV_
package Coefficients_Fx;
	localparam N = 4;
	localparam M = 4;
	localparam COEFF_BIAS = 48;
	localparam logic signed[63:0] Lfr[0:3] = {64'd277509184401256, 64'd277509184401256, 64'd273021858248849, 64'd273021858248849};
	localparam logic signed[63:0] Lfi[0:3] = {64'd16835351421295, - 64'd16835351421295, 64'd6718885687873, - 64'd6718885687873};
	localparam logic signed[63:0] Lbr[0:3] = {64'd277509184401256, 64'd277509184401256, 64'd273021858248849, 64'd273021858248849};
	localparam logic signed[63:0] Lbi[0:3] = {64'd16835351421295, - 64'd16835351421295, 64'd6718885687873, - 64'd6718885687873};
	localparam logic signed[63:0] Wfr[0:3] = {- 64'd9065742652, - 64'd9065742652, 64'd2686576365, 64'd2686576365};
	localparam logic signed[63:0] Wfi[0:3] = {- 64'd399150078, 64'd399150078, 64'd5217631883, - 64'd5217631883};
	localparam logic signed[63:0] Wbr[0:3] = {64'd9065742652, 64'd9065742652, - 64'd2686576365, - 64'd2686576365};
	localparam logic signed[63:0] Wbi[0:3] = {64'd399150078, - 64'd399150078, - 64'd5217631883, 64'd5217631883};
	localparam logic signed[63:0] Ffr[0:3][0:79] = '{
		'{- 64'd26567897873202484, - 64'd3192018314165762, 64'd450274308527086, - 64'd6029254211273, - 64'd28092981743047812, - 64'd2907551920935952, 64'd453015564229319, - 64'd8389181821419, - 64'd29474773437002956, - 64'd2619048706861976, 64'd453979390270136, - 64'd10659844078507, - 64'd30711552191100992, - 64'd2327696536976608, 64'd453205521545409, - 64'd12834845540299, - 64'd31802186785202120, - 64'd2034665046458791, 64'd450739284648358, - 64'd14908308035339, - 64'd32746125427854796, - 64'd1741101669082493, 64'd446631290268612, - 64'd16874880235427, - 64'd33543383700137080, - 64'd1448127846412385, 64'd440937113145429, - 64'd18729745005201, - 64'd34194530651367228, - 64'd1156835427649247, 64'd433716961087251, - 64'd20468624555308, - 64'd34700673144283876, - 64'd868283269066497, 64'd425035334574151, - 64'd22087783433324, - 64'd35063438551524652, - 64'd583494041007436, 64'd414960678458287, - 64'd23584029393878, - 64'd35284955908971984, - 64'd303451249434539, 64'd403565027270315, - 64'd24954712196456, - 64'd35367835634785860, - 64'd29096478041441, 64'd390923645627091, - 64'd26197720385994, - 64'd35315147925703144, 64'd238673144041250, 64'd377114665217978, - 64'd27311476117639, - 64'd35130399944455176, 64'd499007244889776, 64'd362218719823951, - 64'd28294928092948, - 64'd34817511913941216, 64'd751104279690268, 64'd346318579795623, - 64'd29147542680290, - 64'd34380792235101752, 64'd994213365764789, 64'd329498787383581, - 64'd29869293297271, - 64'd33824911746268080, 64'd1227635881523198, 64'd311845294277168, - 64'd30460648137710, - 64'd33154877242132380, 64'd1450726829064212, 64'd293445102666446, - 64'd30922556329883, - 64'd32376004370394872, 64'd1662895961048274, 64'd274385911096659, - 64'd31256432616592, - 64'd31493890023613728, 64'd1863608673339688, 64'd254755766335471, - 64'd31464140650979},
		'{- 64'd26567897873218296, - 64'd3192018314164136, 64'd450274308527077, - 64'd6029254211282, - 64'd28092981743062688, - 64'd2907551920934424, 64'd453015564229310, - 64'd8389181821427, - 64'd29474773437016856, - 64'd2619048706860550, 64'd453979390270128, - 64'd10659844078515, - 64'd30711552191113888, - 64'd2327696536975287, 64'd453205521545401, - 64'd12834845540307, - 64'd31802186785213992, - 64'd2034665046457576, 64'd450739284648350, - 64'd14908308035346, - 64'd32746125427865624, - 64'd1741101669081388, 64'd446631290268605, - 64'd16874880235433, - 64'd33543383700146848, - 64'd1448127846411390, 64'd440937113145422, - 64'd18729745005206, - 64'd34194530651375920, - 64'd1156835427648364, 64'd433716961087244, - 64'd20468624555312, - 64'd34700673144291496, - 64'd868283269065726, 64'd425035334574144, - 64'd22087783433328, - 64'd35063438551531184, - 64'd583494041006778, 64'd414960678458281, - 64'd23584029393881, - 64'd35284955908977440, - 64'd303451249433993, 64'd403565027270309, - 64'd24954712196459, - 64'd35367835634790244, - 64'd29096478041006, 64'd390923645627086, - 64'd26197720385996, - 64'd35315147925706464, 64'd238673144041574, 64'd377114665217974, - 64'd27311476117640, - 64'd35130399944457448, 64'd499007244889991, 64'd362218719823947, - 64'd28294928092949, - 64'd34817511913942448, 64'd751104279690376, 64'd346318579795620, - 64'd29147542680290, - 64'd34380792235101972, 64'd994213365764792, 64'd329498787383578, - 64'd29869293297271, - 64'd33824911746267312, 64'd1227635881523099, 64'd311845294277166, - 64'd30460648137709, - 64'd33154877242130648, 64'd1450726829064013, 64'd293445102666444, - 64'd30922556329881, - 64'd32376004370392208, 64'd1662895961047979, 64'd274385911096657, - 64'd31256432616590, - 64'd31493890023610168, 64'd1863608673339300, 64'd254755766335470, - 64'd31464140650976},
		'{64'd26285687980516512, 64'd3160906636728641, - 64'd428510658795101, 64'd73898504907566, 64'd27799448360287640, 64'd2896044112115250, - 64'd399227411165679, 64'd70470454190196, 64'd29183603555461704, 64'd2642438181955122, - 64'd371072372506860, 64'd67139547471731, 64'd30443710271282672, 64'd2399802534529312, - 64'd344020874801160, 64'd63904994989796, 64'd31585182198078848, 64'd2167851488741114, - 64'd318048071302206, 64'd60765911452485, 64'd32613290423469060, 64'd1946300377598710, - 64'd293128983573209, 64'd57721322938431, 64'd33533164030282976, 64'd1734865907736606, - 64'd269238545963188, 64'd54770173523026, 64'd34349790868434332, 64'd1533266495850688, - 64'd246351647605625, 64'd51911331637084, 64'd35068018489418916, 64'd1341222582904435, - 64'd224443172022907, 64'd49143596164272, 64'd35692555232533728, 64'd1158456926946292, - 64'd203488034418548, 64'd46465702283627, 64'd36227971452329160, 64'd984694875360464, - 64'd183461216737786, 64'd43876327063513, 64'd36678700877212664, 64'd819664617355500, - 64'd164337800575708, 64'd41374094813333, 64'd37049042089520288, 64'd663097417476976, - 64'd146092998010592, 64'd38957582199330, 64'd37343160117760824, 64'd514727830912426, - 64'd128702180438657, 64'd36625323130756, 64'd37565088132116912, 64'd374293901338505, - 64'd112140905484870, 64'd34375813422680, 64'd37718729234658016, 64'd241537342042072, - 64'd96384942062960, 64'd32207515241657, 64'd37807858336081272, 64'd116203701028647, - 64'd81410293656162, 64'd30118861340444, 64'd37836124111148440, - 64'd1957489186539, - 64'd67193219888722, 64'd28108259087881, 64'd37807051025330336, - 64'd113192576427887, - 64'd53710256456519, 64'd26174094300016, 64'd37724041425504024, - 64'd217743667690256, - 64'd40938233483652, 64'd24314734878474},
		'{64'd26285687980563748, 64'd3160906636723780, - 64'd428510658795078, 64'd73898504907594, 64'd27799448360333176, 64'd2896044112110566, - 64'd399227411165656, 64'd70470454190224, 64'd29183603555505572, 64'd2642438181950610, - 64'd371072372506839, 64'd67139547471757, 64'd30443710271324904, 64'd2399802534524968, - 64'd344020874801139, 64'd63904994989821, 64'd31585182198119480, 64'd2167851488736936, - 64'd318048071302186, 64'd60765911452510, 64'd32613290423508120, 64'd1946300377594694, - 64'd293128983573189, 64'd57721322938455, 64'd33533164030320512, 64'd1734865907732748, - 64'd269238545963169, 64'd54770173523048, 64'd34349790868470364, 64'd1533266495846984, - 64'd246351647605607, 64'd51911331637105, 64'd35068018489453484, 64'd1341222582900882, - 64'd224443172022890, 64'd49143596164292, 64'd35692555232566872, 64'd1158456926942886, - 64'd203488034418532, 64'd46465702283647, 64'd36227971452360912, 64'd984694875357202, - 64'd183461216737770, 64'd43876327063532, 64'd36678700877243048, 64'd819664617352380, - 64'd164337800575693, 64'd41374094813351, 64'd37049042089549352, 64'd663097417473992, - 64'd146092998010578, 64'd38957582199348, 64'd37343160117788592, 64'd514727830909575, - 64'd128702180438642, 64'd36625323130773, 64'd37565088132143432, 64'd374293901335783, - 64'd112140905484857, 64'd34375813422696, 64'd37718729234683320, 64'd241537342039476, - 64'd96384942062947, 64'd32207515241672, 64'd37807858336105392, 64'd116203701026173, - 64'd81410293656150, 64'd30118861340458, 64'd37836124111171400, - 64'd1957489188894, - 64'd67193219888710, 64'd28108259087895, 64'd37807051025352184, - 64'd113192576430128, - 64'd53710256456508, 64'd26174094300029, 64'd37724041425524784, - 64'd217743667692384, - 64'd40938233483641, 64'd24314734878486}};
	localparam logic signed[63:0] Ffi[0:3][0:79] = '{
		'{64'd31756730134704588, - 64'd4004151029617032, - 64'd151899963999939, 64'd40876565143546, 64'd29720241846974532, - 64'd4138653638501433, - 64'd122828356908291, 64'd39940025120640, 64'd27621229232884120, - 64'd4254246924888753, - 64'd94002391377932, 64'd38875530251281, 64'd25469143692556908, - 64'd4350955861329947, - 64'd65524916656424, 64'd37690222399226, 64'd23273406383201360, - 64'd4428876116142784, - 64'd37494956323755, 64'd36391525323161, 64'd21043373383899164, - 64'd4488171967007112, - 64'd10007427747382, 64'd34987109766420, 64'd18788301956196616, - 64'd4529074006412982, 64'd16847116112075, 64'd33484858466014, 64'd16517318001154640, - 64'd4551876652704974, 64'd42982722114963, 64'd31892831215079, 64'd14239384806538872, - 64'd4556935480864709, 64'd68318249243579, 64'd30219230109354, 64'd11963273170674172, - 64'd4544664387509117, 64'd92777557552391, 64'd28472365104417, 64'd9697532982177808, - 64'd4515532604854686, 64'd116289673623871, 64'd26660620006160, 64'd7450466327355798, - 64'd4470061578608283, 64'd138788932478523, 64'd24792419012331, 64'd5230102189526454, - 64'd4408821724893831, 64'd160215095977853, 64'd22876193918048, 64'd3044172796956274, - 64'd4332429081412194, 64'd180513447846848, 64'd20920352092900, 64'd900091668485036, - 64'd4241541868060102, 64'd199634865527703, 64'd18933245331719, - 64'd1195066601691070, - 64'd4136856972204280, 64'd217535869158888, 64'd16923139675329, - 64'd3234584786188100, - 64'd4019106373720620, 64'd234178648052799, 64'd14898186291546, - 64'd5212119667186542, - 64'd3889053524766924, 64'd249531065121127, 64'd12866393500509, - 64'd7121716860836634, - 64'd3747489699063430, 64'd263566639769367, 64'd10835600022054, - 64'd8957823811714248, - 64'd3595230325209902, 64'd276264509850467, 64'd8813449516304},
		'{- 64'd31756730134692604, 64'd4004151029615770, 64'd151899963999942, - 64'd40876565143538, - 64'd29720241846961776, 64'd4138653638500091, 64'd122828356908294, - 64'd39940025120632, - 64'd27621229232870648, 64'd4254246924887338, 64'd94002391377935, - 64'd38875530251273, - 64'd25469143692542800, 64'd4350955861328467, 64'd65524916656428, - 64'd37690222399217, - 64'd23273406383186676, 64'd4428876116141246, 64'd37494956323760, - 64'd36391525323152, - 64'd21043373383883972, 64'd4488171967005522, 64'd10007427747387, - 64'd34987109766411, - 64'd18788301956180996, 64'd4529074006411349, - 64'd16847116112070, - 64'd33484858466004, - 64'd16517318001138656, 64'd4551876652703305, - 64'd42982722114958, - 64'd31892831215069, - 64'd14239384806522594, 64'd4556935480863010, - 64'd68318249243573, - 64'd30219230109344, - 64'd11963273170657666, 64'd4544664387507396, - 64'd92777557552385, - 64'd28472365104407, - 64'd9697532982161142, 64'd4515532604852950, - 64'd116289673623865, - 64'd26660620006150, - 64'd7450466327339044, 64'd4470061578606539, - 64'd138788932478516, - 64'd24792419012321, - 64'd5230102189509672, 64'd4408821724892086, - 64'd160215095977846, - 64'd22876193918038, - 64'd3044172796939530, 64'd4332429081410454, - 64'd180513447846841, - 64'd20920352092890, - 64'd900091668468394, 64'd4241541868058373, - 64'd199634865527696, - 64'd18933245331709, 64'd1195066601707554, 64'd4136856972202569, - 64'd217535869158881, - 64'd16923139675319, 64'd3234584786204364, 64'd4019106373718933, - 64'd234178648052792, - 64'd14898186291536, 64'd5212119667202530, 64'd3889053524765268, - 64'd249531065121120, - 64'd12866393500500, 64'd7121716860852294, 64'd3747489699061808, - 64'd263566639769359, - 64'd10835600022045, 64'd8957823811729530, 64'd3595230325208320, - 64'd276264509850460, - 64'd8813449516294},
		'{- 64'd96486490782400608, 64'd7119135065273385, - 64'd687651241321332, 64'd50639004070964, - 64'd92961409153791744, 64'd6980788409576997, - 64'd677228704635829, 64'd50882216123342, - 64'd89506057168197776, 64'd6840274170944421, - 64'd666420173225727, 64'd51036295630137, - 64'd86121434450844496, 64'd6697926143192068, - 64'd655264169756044, 64'd51106238230416, - 64'd82808377966609312, 64'd6554061261464093, - 64'd643797471165597, 64'd51096870684820, - 64'd79567570318762688, 64'd6408980123576888, - 64'd632055156827496, 64'd51012853666916, - 64'd76399547788646352, 64'd6262967504860670, - 64'd620070656386110, 64'd50858684635437, - 64'd73304708119635456, 64'd6116292866121464, - 64'd607875797219092, 64'd50638700778427, - 64'd70283318048911624, 64'd5969210854379020, - 64'd595500851476554, 64'd50357082020754, - 64'd67335520590738840, 64'd5821961796067011, - 64'd582974582652960, 64'd50017854086856, - 64'd64461342075083248, 64'd5674772182411308, - 64'd570324291650575, 64'd49624891610959, - 64'd61660698945552744, 64'd5527855146730314, - 64'd557575862296453, 64'd49181921287432, - 64'd58933404320754288, 64'd5381410933428235, - 64'd544753806278019, 64'd48692525054269, - 64'd56279174323273712, 64'd5235627358477770, - 64'd531881307465164, 64'd48160143303088, - 64'd53697634180579488, 64'd5090680261213204, - 64'd518980265589570, 64'd47588078109359, - 64'd51188324102235200, 64'd4946733947278150, - 64'd506071339254650, 64'd46979496476934, - 64'd48750704937877416, 64'd4803941622594292, - 64'd493173988252031, 64'd46337433591244, - 64'd46384163620477680, 64'd4662445818238601, - 64'd480306515162914, 64'd45664796075895, - 64'd44088018399458320, 64'd4522378806136374, - 64'd467486106225012, 64'd44964365247652, - 64'd41861523868273272, 64'd4383863005496490, - 64'd454728871447932, 64'd44238800365119},
		'{64'd96486490782388784, - 64'd7119135065272138, 64'd687651241321330, - 64'd50639004070972, 64'd92961409153779168, - 64'd6980788409575672, 64'd677228704635826, - 64'd50882216123350, 64'd89506057168184464, - 64'd6840274170943023, 64'd666420173225724, - 64'd51036295630145, 64'd86121434450830544, - 64'd6697926143190605, 64'd655264169756040, - 64'd51106238230425, 64'd82808377966594784, - 64'd6554061261462569, 64'd643797471165593, - 64'd51096870684829, 64'd79567570318747616, - 64'd6408980123575310, 64'd632055156827491, - 64'd51012853666926, 64'd76399547788630800, - 64'd6262967504859045, 64'd620070656386106, - 64'd50858684635447, 64'd73304708119619472, - 64'd6116292866119796, 64'd607875797219087, - 64'd50638700778437, 64'd70283318048895248, - 64'd5969210854377313, 64'd595500851476548, - 64'd50357082020764, 64'd67335520590722136, - 64'd5821961796065270, 64'd582974582652954, - 64'd50017854086866, 64'd64461342075066256, - 64'd5674772182409537, 64'd570324291650569, - 64'd49624891610970, 64'd61660698945535520, - 64'd5527855146728520, 64'd557575862296446, - 64'd49181921287443, 64'd58933404320736848, - 64'd5381410933426420, 64'd544753806278013, - 64'd48692525054280, 64'd56279174323256096, - 64'd5235627358475938, 64'd531881307465158, - 64'd48160143303099, 64'd53697634180561744, - 64'd5090680261211360, 64'd518980265589563, - 64'd47588078109370, 64'd51188324102217360, - 64'd4946733947276296, 64'd506071339254643, - 64'd46979496476945, 64'd48750704937859504, - 64'd4803941622592431, 64'd493173988252024, - 64'd46337433591255, 64'd46384163620459736, - 64'd4662445818236737, 64'd480306515162907, - 64'd45664796075906, 64'd44088018399440360, - 64'd4522378806134510, 64'd467486106225005, - 64'd44964365247663, 64'd41861523868255320, - 64'd4383863005494629, 64'd454728871447925, - 64'd44238800365130}};
	localparam logic signed[63:0] Fbr[0:3][0:79] = '{
		'{64'd26567897873202484, - 64'd3192018314165762, - 64'd450274308527086, - 64'd6029254211273, 64'd28092981743047812, - 64'd2907551920935952, - 64'd453015564229319, - 64'd8389181821419, 64'd29474773437002956, - 64'd2619048706861976, - 64'd453979390270136, - 64'd10659844078507, 64'd30711552191100992, - 64'd2327696536976608, - 64'd453205521545409, - 64'd12834845540299, 64'd31802186785202120, - 64'd2034665046458791, - 64'd450739284648358, - 64'd14908308035339, 64'd32746125427854796, - 64'd1741101669082493, - 64'd446631290268612, - 64'd16874880235427, 64'd33543383700137080, - 64'd1448127846412385, - 64'd440937113145429, - 64'd18729745005201, 64'd34194530651367228, - 64'd1156835427649247, - 64'd433716961087251, - 64'd20468624555308, 64'd34700673144283876, - 64'd868283269066497, - 64'd425035334574151, - 64'd22087783433324, 64'd35063438551524652, - 64'd583494041007436, - 64'd414960678458287, - 64'd23584029393878, 64'd35284955908971984, - 64'd303451249434539, - 64'd403565027270315, - 64'd24954712196456, 64'd35367835634785860, - 64'd29096478041441, - 64'd390923645627091, - 64'd26197720385994, 64'd35315147925703144, 64'd238673144041250, - 64'd377114665217978, - 64'd27311476117639, 64'd35130399944455176, 64'd499007244889776, - 64'd362218719823951, - 64'd28294928092948, 64'd34817511913941216, 64'd751104279690268, - 64'd346318579795623, - 64'd29147542680290, 64'd34380792235101752, 64'd994213365764789, - 64'd329498787383581, - 64'd29869293297271, 64'd33824911746268080, 64'd1227635881523198, - 64'd311845294277168, - 64'd30460648137710, 64'd33154877242132380, 64'd1450726829064212, - 64'd293445102666446, - 64'd30922556329883, 64'd32376004370394872, 64'd1662895961048274, - 64'd274385911096659, - 64'd31256432616592, 64'd31493890023613728, 64'd1863608673339688, - 64'd254755766335471, - 64'd31464140650979},
		'{64'd26567897873218296, - 64'd3192018314164136, - 64'd450274308527077, - 64'd6029254211282, 64'd28092981743062688, - 64'd2907551920934424, - 64'd453015564229310, - 64'd8389181821427, 64'd29474773437016856, - 64'd2619048706860550, - 64'd453979390270128, - 64'd10659844078515, 64'd30711552191113888, - 64'd2327696536975287, - 64'd453205521545401, - 64'd12834845540307, 64'd31802186785213992, - 64'd2034665046457576, - 64'd450739284648350, - 64'd14908308035346, 64'd32746125427865624, - 64'd1741101669081388, - 64'd446631290268605, - 64'd16874880235433, 64'd33543383700146848, - 64'd1448127846411390, - 64'd440937113145422, - 64'd18729745005206, 64'd34194530651375920, - 64'd1156835427648364, - 64'd433716961087244, - 64'd20468624555312, 64'd34700673144291496, - 64'd868283269065726, - 64'd425035334574144, - 64'd22087783433328, 64'd35063438551531184, - 64'd583494041006778, - 64'd414960678458281, - 64'd23584029393881, 64'd35284955908977440, - 64'd303451249433993, - 64'd403565027270309, - 64'd24954712196459, 64'd35367835634790244, - 64'd29096478041006, - 64'd390923645627086, - 64'd26197720385996, 64'd35315147925706464, 64'd238673144041574, - 64'd377114665217974, - 64'd27311476117640, 64'd35130399944457448, 64'd499007244889991, - 64'd362218719823947, - 64'd28294928092949, 64'd34817511913942448, 64'd751104279690376, - 64'd346318579795620, - 64'd29147542680290, 64'd34380792235101972, 64'd994213365764792, - 64'd329498787383578, - 64'd29869293297271, 64'd33824911746267312, 64'd1227635881523099, - 64'd311845294277166, - 64'd30460648137709, 64'd33154877242130648, 64'd1450726829064013, - 64'd293445102666444, - 64'd30922556329881, 64'd32376004370392208, 64'd1662895961047979, - 64'd274385911096657, - 64'd31256432616590, 64'd31493890023610168, 64'd1863608673339300, - 64'd254755766335470, - 64'd31464140650976},
		'{- 64'd26285687980516512, 64'd3160906636728641, 64'd428510658795101, 64'd73898504907566, - 64'd27799448360287640, 64'd2896044112115250, 64'd399227411165679, 64'd70470454190196, - 64'd29183603555461704, 64'd2642438181955122, 64'd371072372506860, 64'd67139547471731, - 64'd30443710271282672, 64'd2399802534529312, 64'd344020874801160, 64'd63904994989796, - 64'd31585182198078848, 64'd2167851488741114, 64'd318048071302206, 64'd60765911452485, - 64'd32613290423469060, 64'd1946300377598710, 64'd293128983573209, 64'd57721322938431, - 64'd33533164030282976, 64'd1734865907736606, 64'd269238545963188, 64'd54770173523026, - 64'd34349790868434332, 64'd1533266495850688, 64'd246351647605625, 64'd51911331637084, - 64'd35068018489418916, 64'd1341222582904435, 64'd224443172022907, 64'd49143596164272, - 64'd35692555232533728, 64'd1158456926946292, 64'd203488034418548, 64'd46465702283627, - 64'd36227971452329160, 64'd984694875360464, 64'd183461216737786, 64'd43876327063513, - 64'd36678700877212664, 64'd819664617355500, 64'd164337800575708, 64'd41374094813333, - 64'd37049042089520288, 64'd663097417476976, 64'd146092998010592, 64'd38957582199330, - 64'd37343160117760824, 64'd514727830912426, 64'd128702180438657, 64'd36625323130756, - 64'd37565088132116912, 64'd374293901338505, 64'd112140905484870, 64'd34375813422680, - 64'd37718729234658016, 64'd241537342042072, 64'd96384942062960, 64'd32207515241657, - 64'd37807858336081272, 64'd116203701028647, 64'd81410293656162, 64'd30118861340444, - 64'd37836124111148440, - 64'd1957489186539, 64'd67193219888722, 64'd28108259087881, - 64'd37807051025330336, - 64'd113192576427887, 64'd53710256456519, 64'd26174094300016, - 64'd37724041425504024, - 64'd217743667690256, 64'd40938233483652, 64'd24314734878474},
		'{- 64'd26285687980563748, 64'd3160906636723780, 64'd428510658795078, 64'd73898504907594, - 64'd27799448360333176, 64'd2896044112110566, 64'd399227411165656, 64'd70470454190224, - 64'd29183603555505572, 64'd2642438181950610, 64'd371072372506839, 64'd67139547471757, - 64'd30443710271324904, 64'd2399802534524968, 64'd344020874801139, 64'd63904994989821, - 64'd31585182198119480, 64'd2167851488736936, 64'd318048071302186, 64'd60765911452510, - 64'd32613290423508120, 64'd1946300377594694, 64'd293128983573189, 64'd57721322938455, - 64'd33533164030320512, 64'd1734865907732748, 64'd269238545963169, 64'd54770173523048, - 64'd34349790868470364, 64'd1533266495846984, 64'd246351647605607, 64'd51911331637105, - 64'd35068018489453484, 64'd1341222582900882, 64'd224443172022890, 64'd49143596164292, - 64'd35692555232566872, 64'd1158456926942886, 64'd203488034418532, 64'd46465702283647, - 64'd36227971452360912, 64'd984694875357202, 64'd183461216737770, 64'd43876327063532, - 64'd36678700877243048, 64'd819664617352380, 64'd164337800575693, 64'd41374094813351, - 64'd37049042089549352, 64'd663097417473992, 64'd146092998010578, 64'd38957582199348, - 64'd37343160117788592, 64'd514727830909575, 64'd128702180438642, 64'd36625323130773, - 64'd37565088132143432, 64'd374293901335783, 64'd112140905484857, 64'd34375813422696, - 64'd37718729234683320, 64'd241537342039476, 64'd96384942062947, 64'd32207515241672, - 64'd37807858336105392, 64'd116203701026173, 64'd81410293656150, 64'd30118861340458, - 64'd37836124111171400, - 64'd1957489188894, 64'd67193219888710, 64'd28108259087895, - 64'd37807051025352184, - 64'd113192576430128, 64'd53710256456508, 64'd26174094300029, - 64'd37724041425524784, - 64'd217743667692384, 64'd40938233483641, 64'd24314734878486}};
	localparam logic signed[63:0] Fbi[0:3][0:79] = '{
		'{- 64'd31756730134704588, - 64'd4004151029617032, 64'd151899963999939, 64'd40876565143546, - 64'd29720241846974532, - 64'd4138653638501433, 64'd122828356908291, 64'd39940025120640, - 64'd27621229232884120, - 64'd4254246924888753, 64'd94002391377932, 64'd38875530251281, - 64'd25469143692556908, - 64'd4350955861329947, 64'd65524916656424, 64'd37690222399226, - 64'd23273406383201360, - 64'd4428876116142784, 64'd37494956323755, 64'd36391525323161, - 64'd21043373383899164, - 64'd4488171967007112, 64'd10007427747382, 64'd34987109766420, - 64'd18788301956196616, - 64'd4529074006412982, - 64'd16847116112075, 64'd33484858466014, - 64'd16517318001154640, - 64'd4551876652704974, - 64'd42982722114963, 64'd31892831215079, - 64'd14239384806538872, - 64'd4556935480864709, - 64'd68318249243579, 64'd30219230109354, - 64'd11963273170674172, - 64'd4544664387509117, - 64'd92777557552391, 64'd28472365104417, - 64'd9697532982177808, - 64'd4515532604854686, - 64'd116289673623871, 64'd26660620006160, - 64'd7450466327355798, - 64'd4470061578608283, - 64'd138788932478523, 64'd24792419012331, - 64'd5230102189526454, - 64'd4408821724893831, - 64'd160215095977853, 64'd22876193918048, - 64'd3044172796956274, - 64'd4332429081412194, - 64'd180513447846848, 64'd20920352092900, - 64'd900091668485036, - 64'd4241541868060102, - 64'd199634865527703, 64'd18933245331719, 64'd1195066601691070, - 64'd4136856972204280, - 64'd217535869158888, 64'd16923139675329, 64'd3234584786188100, - 64'd4019106373720620, - 64'd234178648052799, 64'd14898186291546, 64'd5212119667186542, - 64'd3889053524766924, - 64'd249531065121127, 64'd12866393500509, 64'd7121716860836634, - 64'd3747489699063430, - 64'd263566639769367, 64'd10835600022054, 64'd8957823811714248, - 64'd3595230325209902, - 64'd276264509850467, 64'd8813449516304},
		'{64'd31756730134692604, 64'd4004151029615770, - 64'd151899963999942, - 64'd40876565143538, 64'd29720241846961776, 64'd4138653638500091, - 64'd122828356908294, - 64'd39940025120632, 64'd27621229232870648, 64'd4254246924887338, - 64'd94002391377935, - 64'd38875530251273, 64'd25469143692542800, 64'd4350955861328467, - 64'd65524916656428, - 64'd37690222399217, 64'd23273406383186676, 64'd4428876116141246, - 64'd37494956323760, - 64'd36391525323152, 64'd21043373383883972, 64'd4488171967005522, - 64'd10007427747387, - 64'd34987109766411, 64'd18788301956180996, 64'd4529074006411349, 64'd16847116112070, - 64'd33484858466004, 64'd16517318001138656, 64'd4551876652703305, 64'd42982722114958, - 64'd31892831215069, 64'd14239384806522594, 64'd4556935480863010, 64'd68318249243573, - 64'd30219230109344, 64'd11963273170657666, 64'd4544664387507396, 64'd92777557552385, - 64'd28472365104407, 64'd9697532982161142, 64'd4515532604852950, 64'd116289673623865, - 64'd26660620006150, 64'd7450466327339044, 64'd4470061578606539, 64'd138788932478516, - 64'd24792419012321, 64'd5230102189509672, 64'd4408821724892086, 64'd160215095977846, - 64'd22876193918038, 64'd3044172796939530, 64'd4332429081410454, 64'd180513447846841, - 64'd20920352092890, 64'd900091668468394, 64'd4241541868058373, 64'd199634865527696, - 64'd18933245331709, - 64'd1195066601707554, 64'd4136856972202569, 64'd217535869158881, - 64'd16923139675319, - 64'd3234584786204364, 64'd4019106373718933, 64'd234178648052792, - 64'd14898186291536, - 64'd5212119667202530, 64'd3889053524765268, 64'd249531065121120, - 64'd12866393500500, - 64'd7121716860852294, 64'd3747489699061808, 64'd263566639769359, - 64'd10835600022045, - 64'd8957823811729530, 64'd3595230325208320, 64'd276264509850460, - 64'd8813449516294},
		'{64'd96486490782400608, 64'd7119135065273385, 64'd687651241321332, 64'd50639004070964, 64'd92961409153791744, 64'd6980788409576997, 64'd677228704635829, 64'd50882216123342, 64'd89506057168197776, 64'd6840274170944421, 64'd666420173225727, 64'd51036295630137, 64'd86121434450844496, 64'd6697926143192068, 64'd655264169756044, 64'd51106238230416, 64'd82808377966609312, 64'd6554061261464093, 64'd643797471165597, 64'd51096870684820, 64'd79567570318762688, 64'd6408980123576888, 64'd632055156827496, 64'd51012853666916, 64'd76399547788646352, 64'd6262967504860670, 64'd620070656386110, 64'd50858684635437, 64'd73304708119635456, 64'd6116292866121464, 64'd607875797219092, 64'd50638700778427, 64'd70283318048911624, 64'd5969210854379020, 64'd595500851476554, 64'd50357082020754, 64'd67335520590738840, 64'd5821961796067011, 64'd582974582652960, 64'd50017854086856, 64'd64461342075083248, 64'd5674772182411308, 64'd570324291650575, 64'd49624891610959, 64'd61660698945552744, 64'd5527855146730314, 64'd557575862296453, 64'd49181921287432, 64'd58933404320754288, 64'd5381410933428235, 64'd544753806278019, 64'd48692525054269, 64'd56279174323273712, 64'd5235627358477770, 64'd531881307465164, 64'd48160143303088, 64'd53697634180579488, 64'd5090680261213204, 64'd518980265589570, 64'd47588078109359, 64'd51188324102235200, 64'd4946733947278150, 64'd506071339254650, 64'd46979496476934, 64'd48750704937877416, 64'd4803941622594292, 64'd493173988252031, 64'd46337433591244, 64'd46384163620477680, 64'd4662445818238601, 64'd480306515162914, 64'd45664796075895, 64'd44088018399458320, 64'd4522378806136374, 64'd467486106225012, 64'd44964365247652, 64'd41861523868273272, 64'd4383863005496490, 64'd454728871447932, 64'd44238800365119},
		'{- 64'd96486490782388784, - 64'd7119135065272138, - 64'd687651241321330, - 64'd50639004070972, - 64'd92961409153779168, - 64'd6980788409575672, - 64'd677228704635826, - 64'd50882216123350, - 64'd89506057168184464, - 64'd6840274170943023, - 64'd666420173225724, - 64'd51036295630145, - 64'd86121434450830544, - 64'd6697926143190605, - 64'd655264169756040, - 64'd51106238230425, - 64'd82808377966594784, - 64'd6554061261462569, - 64'd643797471165593, - 64'd51096870684829, - 64'd79567570318747616, - 64'd6408980123575310, - 64'd632055156827491, - 64'd51012853666926, - 64'd76399547788630800, - 64'd6262967504859045, - 64'd620070656386106, - 64'd50858684635447, - 64'd73304708119619472, - 64'd6116292866119796, - 64'd607875797219087, - 64'd50638700778437, - 64'd70283318048895248, - 64'd5969210854377313, - 64'd595500851476548, - 64'd50357082020764, - 64'd67335520590722136, - 64'd5821961796065270, - 64'd582974582652954, - 64'd50017854086866, - 64'd64461342075066256, - 64'd5674772182409537, - 64'd570324291650569, - 64'd49624891610970, - 64'd61660698945535520, - 64'd5527855146728520, - 64'd557575862296446, - 64'd49181921287443, - 64'd58933404320736848, - 64'd5381410933426420, - 64'd544753806278013, - 64'd48692525054280, - 64'd56279174323256096, - 64'd5235627358475938, - 64'd531881307465158, - 64'd48160143303099, - 64'd53697634180561744, - 64'd5090680261211360, - 64'd518980265589563, - 64'd47588078109370, - 64'd51188324102217360, - 64'd4946733947276296, - 64'd506071339254643, - 64'd46979496476945, - 64'd48750704937859504, - 64'd4803941622592431, - 64'd493173988252024, - 64'd46337433591255, - 64'd46384163620459736, - 64'd4662445818236737, - 64'd480306515162907, - 64'd45664796075906, - 64'd44088018399440360, - 64'd4522378806134510, - 64'd467486106225005, - 64'd44964365247663, - 64'd41861523868255320, - 64'd4383863005494629, - 64'd454728871447925, - 64'd44238800365130}};
	localparam logic signed[63:0] hf[0:1199] = {64'd5880330321920, - 64'd9331200000, - 64'd12121982976, 64'd37615036, 64'd5871003762688, - 64'd27963885568, - 64'd12043516928, 64'd112520208, 64'd5852380528640, - 64'd46507737088, - 64'd11887098880, 64'd186471232, 64'd5824520388608, - 64'd64904146944, - 64'd11653682176, 64'd258876112, 64'd5787510374400, - 64'd83095248896, - 64'd11344629760, 64'd329181408, 64'd5741467926528, - 64'd101024178176, - 64'd10961692672, 64'd396872800, 64'd5686538797056, - 64'd118635307008, - 64'd10506989568, 64'd461475424, 64'd5622894428160, - 64'd135874502656, - 64'd9982984192, 64'd522554208, 64'd5550734573568, - 64'd152689360896, - 64'd9392459776, 64'd579713856, 64'd5470283628544, - 64'd169029353472, - 64'd8738495488, 64'd632598976, 64'd5381791678464, - 64'd184846123008, - 64'd8024443392, 64'd680893760, 64'd5285531877376, - 64'd200093564928, - 64'd7253902336, 64'd724321536, 64'd5181799923712, - 64'd214728081408, - 64'd6430694400, 64'd762644672, 64'd5070912487424, - 64'd228708646912, - 64'd5558839296, 64'd795663808, 64'd4953206685696, - 64'd241997037568, - 64'd4642529792, 64'd823217088, 64'd4829036412928, - 64'd254557880320, - 64'd3686106112, 64'd845179392, 64'd4698774962176, - 64'd266358784000, - 64'd2694032896, 64'd861461696, 64'd4562809257984, - 64'd277370437632, - 64'd1670873728, 64'd872009664, 64'd4421540380672, - 64'd287566626816, - 64'd621268032, 64'd876802624, 64'd4275381993472, - 64'd296924446720, 64'd450092960, 64'd875852672, 64'd4124758769664, - 64'd305424171008, 64'd1538488960, 64'd869203008, 64'd3970103508992, - 64'd313049317376, 64'd2639193088, 64'd856926848, 64'd3811857137664, - 64'd319786811392, 64'd3747492864, 64'd839125696, 64'd3650466086912, - 64'd325626822656, 64'd4858712576, 64'd815928384, 64'd3486380982272, - 64'd330562732032, 64'd5968231424, 64'd787488832, 64'd3320054546432, - 64'd334591328256, 64'd7071505408, 64'd753985088, 64'd3151940812800, - 64'd337712480256, 64'd8164083712, 64'd715617280, 64'd2982492766208, - 64'd339929333760, 64'd9241626624, 64'd672606272, 64'd2812161032192, - 64'd341248049152, 64'd10299923456, 64'd625191680, 64'd2641392828416, - 64'd341677899776, 64'd11334905856, 64'd573630336, 64'd2470629343232, - 64'd341231042560, 64'd12342664192, 64'd518194528, 64'd2300305211392, - 64'd339922550784, 64'd13319460864, 64'd459170304, 64'd2130847334400, - 64'd337770184704, 64'd14261741568, 64'd396855712, 64'd1962672390144, - 64'd334794358784, 64'd15166146560, 64'd331559072, 64'd1796186439680, - 64'd331017977856, 64'd16029522944, 64'd263597264, 64'd1631783616512, - 64'd326466371584, 64'd16848930816, 64'd193294128, 64'd1469844684800, - 64'd321167097856, 64'd17621653504, 64'd120978672, 64'd1310736252928, - 64'd315149746176, 64'd18345203712, 64'd46983556, 64'd1154809462784, - 64'd308446003200, 64'd19017326592, - 64'd28356576, 64'd1002399203328, - 64'd301089226752, 64'd19636006912, - 64'd104706624, 64'd853823324160, - 64'd293114478592, 64'd20199477248, - 64'd181732544, 64'd709381718016, - 64'd284558295040, 64'd20706205696, - 64'd259102800, 64'd569355730944, - 64'd275458523136, 64'd21154916352, - 64'd336489792, 64'd434007375872, - 64'd265854238720, 64'd21544572928, - 64'd413571200, 64'd303579004928, - 64'd255785402368, 64'd21874386944, - 64'd490031264, 64'd178292686848, - 64'd245292875776, 64'd22143815680, - 64'd565561984, 64'd58349928448, - 64'd234418176000, 64'd22352556032, - 64'd639864384, - 64'd56068689920, - 64'd223203344384, 64'd22500540416, - 64'd712649344, - 64'd164803657728, - 64'd211690684416, 64'd22587938816, - 64'd783638912, - 64'd267716722688, - 64'd199922761728, 64'd22615146496, - 64'd852567168, - 64'd364690866176, - 64'd187942109184, 64'd22582779904, - 64'd919180992, - 64'd455630323712, - 64'd175791144960, 64'd22491672576, - 64'd983240768, - 64'd540460515328, - 64'd163512008704, 64'd22342860800, - 64'd1044521472, - 64'd619127832576, - 64'd151146397696, 64'd22137585664, - 64'd1102812928, - 64'd691599245312, - 64'd138735403008, 64'd21877274624, - 64'd1157920384, - 64'd757862301696, - 64'd126319476736, 64'd21563535360, - 64'd1209665408, - 64'd817924407296, - 64'd113938153472, 64'd21198149632, - 64'd1257885696, - 64'd871812562944, - 64'd101630058496, 64'd20783056896, - 64'd1302435840, - 64'd919572840448, - 64'd89432686592, 64'd20320348160, - 64'd1343187328, - 64'd961269661696, - 64'd77382361088, 64'd19812251648, - 64'd1380028928, - 64'd996985405440, - 64'd65514090496, 64'd19261124608, - 64'd1412866432, - 64'd1026819620864, - 64'd53861486592, 64'd18669438976, - 64'd1441623168, - 64'd1050888110080, - 64'd42456657920, 64'd18039771136, - 64'd1466239488, - 64'd1069322600448, - 64'd31330148352, 64'd17374785536, - 64'd1486672896, - 64'd1082269433856, - 64'd20510838784, 64'd16677234688, - 64'd1502897792, - 64'd1089889107968, - 64'd10025896960, 64'd15949931520, - 64'd1514905216, - 64'd1092355227648, 64'd99294480, 64'd15195747328, - 64'd1522702848, - 64'd1089853652992, 64'd9841181696, 64'd14417598464, - 64'd1526313984, - 64'd1082581450752, 64'd19178088448, 64'd13618429952, - 64'd1525777664, - 64'd1070746304512, 64'd28090251264, 64'd12801209344, - 64'd1521148160, - 64'd1054564941824, 64'd36559847424, 64'd11968911360, - 64'd1512493952, - 64'd1034262806528, 64'd44571013120, 64'd11124508672, - 64'd1499897856, - 64'd1010072616960, 64'd52109860864, 64'd10270958592, - 64'd1483456128, - 64'd982233645056, 64'd59164479488, 64'd9411194880, - 64'd1463277440, - 64'd950990536704, 64'd65724940288, 64'd8548114432, - 64'd1439482880, - 64'd916592394240, 64'd71783268352, 64'd7684571136, - 64'd1412204416, - 64'd879291924480, 64'd77333463040, 64'd6823361024, - 64'd1381585280, - 64'd839344324608, 64'd82371428352, 64'd5967217664, - 64'd1347777792, - 64'd797006233600, 64'd86894968832, 64'd5118800896, - 64'd1310943872, - 64'd752535142400, 64'd90903748608, 64'd4280687872, - 64'd1271253504, - 64'd706188083200, 64'd94399275008, 64'd3455368448, - 64'd1228883712, - 64'd658220908544, 64'd97384783872, 64'd2645234176, - 64'd1184018688, - 64'd608887504896, 64'd99865255936, 64'd1852573824, - 64'd1136848000, - 64'd558438744064, 64'd101847326720, 64'd1079566336, - 64'd1087566080, - 64'd507121893376, 64'd103339220992, 64'd328275104, - 64'd1036371520, - 64'd455179632640, 64'd104350679040, - 64'd399356832, - 64'd983466112, - 64'd402849431552, 64'd104892923904, - 64'd1101511680, - 64'd929053952, - 64'd350362861568, 64'd104978538496, - 64'd1776500480, - 64'd873340736, - 64'd297944743936, 64'd104621391872, - 64'd2422767104, - 64'd816532992, - 64'd245812789248, 64'd103836614656, - 64'd3038890496, - 64'd758836928, - 64'd194176761856, 64'd102640427008, - 64'd3623587072, - 64'd700458176, - 64'd143238103040, 64'd101050114048, - 64'd4175712512, - 64'd641600704, - 64'd93189341184, 64'd99083935744, - 64'd4694262784, - 64'd582466112, - 64'd44213682176, 64'd96760987648, - 64'd5178375168, - 64'd523253056, 64'd3515442688, 64'd94101176320, - 64'd5627326976, - 64'd464156384, 64'd49834721280, 64'd91125080064, - 64'd6040537088, - 64'd405366656, 64'd94591270912, 64'd87853858816, - 64'd6417562624, - 64'd347069472, 64'd137642950656, 64'd84309204992, - 64'd6758099456, - 64'd289444800, 64'd178858524672, 64'd80513187840, - 64'd7061979136, - 64'd232666592, 64'd218117931008, 64'd76488237056, - 64'd7329165824, - 64'd176902112, 64'd255312314368, 64'd72256970752, - 64'd7559755264, - 64'd122311512, 64'd290344239104, 64'd67842166784, - 64'd7753970176, - 64'd69047432, 64'd323127640064, 64'd63266664448, - 64'd7912156160, - 64'd17254548, 64'd353587888128, 64'd58553266176, - 64'd8034778112, 64'd32930780, 64'd381661642752, 64'd53724651520, - 64'd8122417152, 64'd81380816, 64'd407297032192, 64'd48803319808, - 64'd8175762432, 64'd127976752, 64'd430453161984, 64'd43811487744, - 64'd8195609600, 64'd172608928, 64'd451100344320, 64'd38771027968, - 64'd8182854144, 64'd215177056, 64'd469219639296, 64'd33703397376, - 64'd8138483712, 64'd255590368, 64'd484802691072, 64'd28629559296, - 64'd8063577088, 64'd293767776, 64'd497851531264, 64'd23569926144, - 64'd7959292416, 64'd329637856, 64'd508378251264, 64'd18544300032, - 64'd7826866176, 64'd363139040, 64'd516404641792, 64'd13571805184, - 64'd7667602432, 64'd394219488, 64'd521961930752, 64'd8670844928, - 64'd7482871296, 64'd422837184, 64'd525090324480, 64'd3859045632, - 64'd7274096640, 64'd448959712, 64'd525838614528, - 64'd846788480, - 64'd7042754560, 64'd472564352, 64'd524263817216, - 64'd5430713856, - 64'd6790364160, 64'd493637728, 64'd520430714880, - 64'd9877687296, - 64'd6518481408, 64'd512175872, 64'd514411298816, - 64'd14173598720, - 64'd6228693504, 64'd528183840, 64'd506284474368, - 64'd18305296384, - 64'd5922609664, 64'd541675520, 64'd496135405568, - 64'd22260619264, - 64'd5601858560, 64'd552673600, 64'd484055089152, - 64'd26028408832, - 64'd5268078080, 64'd561208832, 64'd470139928576, - 64'd29598525440, - 64'd4922912768, 64'd567320192, 64'd454491045888, - 64'd32961867776, - 64'd4568003584, 64'd571054272, 64'd437213855744, - 64'd36110372864, - 64'd4204985344, 64'd572465024, 64'd418417639424, - 64'd39037022208, - 64'd3835479296, 64'd571613376, 64'd398214823936, - 64'd41735839744, - 64'd3461087744, 64'd568566912, 64'd376720621568, - 64'd44201889792, - 64'd3083388160, 64'd563399296, 64'd354052407296, - 64'd46431268864, - 64'd2703929344, 64'd556190080, 64'd330329292800, - 64'd48421093376, - 64'd2324225024, 64'd547024064, 64'd305671569408, - 64'd50169475072, - 64'd1945749504, 64'd535990976, 64'd280200216576, - 64'd51675516928, - 64'd1569933696, 64'd523185088, 64'd254036443136, - 64'd52939288576, - 64'd1198160256, 64'd508704608, 64'd227301163008, - 64'd53961793536, - 64'd831760256, 64'd492651296, 64'd200114569216, - 64'd54744944640, - 64'd472009056, 64'd475130048, 64'd172595675136, - 64'd55291535360, - 64'd120123344, 64'd456248384, 64'd144861888512, - 64'd55605202944, 64'd222742160, 64'd436116000, 64'd117028585472, - 64'd55690399744, 64'd555497280, 64'd414844320, 64'd89208733696, - 64'd55552348160, 64'd877118976, 64'd392546016, 64'd61512495104, - 64'd55196999680, 64'd1186653184, 64'd369334656, 64'd34046879744, - 64'd54631010304, 64'd1483216768, 64'd345324096, 64'd6915413504, - 64'd53861675008, 64'd1765999360, 64'd320628256, - 64'd19782180864, - 64'd52896890880, 64'd2034263808, 64'd295360544, - 64'd45950271488, - 64'd51745124352, 64'd2287347712, 64'd269633472, - 64'd71497596928, - 64'd50415345664, 64'd2524663808, 64'd243558400, - 64'd96337477632, - 64'd48916996096, 64'd2745700096, 64'd217244960, - 64'd120388091904, - 64'd47259926528, 64'd2950020096, 64'd190800800, - 64'd143572615168, - 64'd45454368768, 64'd3137262336, 64'd164331248, - 64'd165819432960, - 64'd43510865920, 64'd3307140096, 64'd137938944, - 64'd187062255616, - 64'd41440239616, 64'd3459440128, 64'd111723488, - 64'd207240282112, - 64'd39253532672, 64'd3594022400, 64'd85781248, - 64'd226298265600, - 64'd36961959936, 64'd3710817792, 64'd60205020, - 64'd244186611712, - 64'd34576879616, 64'd3809826816, 64'd35083764, - 64'd260861427712, - 64'd32109721600, 64'd3891118848, 64'd10502396, - 64'd276284538880, - 64'd29571948544, 64'd3954828288, - 64'd13458433, - 64'd290423472128, - 64'd26975027200, 64'd4001154304, - 64'd36722532, - 64'd303251554304, - 64'd24330364928, 64'd4030357248, - 64'd59218340, - 64'd314747748352, - 64'd21649278976, 64'd4042756096, - 64'd80879072, - 64'd324896587776, - 64'd18942945280, 64'd4038726400, - 64'd101642872, - 64'd333688274944, - 64'd16222372864, 64'd4018696960, - 64'd121452864, - 64'd341118353408, - 64'd13498356736, 64'd3983147776, - 64'd140257312, - 64'd347187773440, - 64'd10781442048, 64'd3932604928, - 64'd158009632, - 64'd351902662656, - 64'd8081892864, 64'd3867639552, - 64'd174668432, - 64'd355274194944, - 64'd5409659904, 64'd3788863488, - 64'd190197584, - 64'd357318459392, - 64'd2774347008, 64'd3696925696, - 64'd204566176, - 64'd358056230912, - 64'd185187008, 64'd3592510208, - 64'd217748528, - 64'd357512806400, 64'd2348986880, 64'd3476330752, - 64'd229724128, - 64'd355717775360, 64'd4819764224, 64'd3349128448, - 64'd240477616, - 64'd352704888832, 64'd7219179520, 64'd3211668736, - 64'd249998672, - 64'd348511731712, 64'd9539730432, 64'd3064736512, - 64'd258281952, - 64'd343179460608, 64'd11774398464, 64'd2909133824, - 64'd265326992, - 64'd336752738304, 64'd13916656640, 64'd2745675776, - 64'd271138016, - 64'd329279209472, 64'd15960493056, 64'd2575187456, - 64'd275723936, - 64'd320809533440, 64'd17900410880, 64'd2398499840, - 64'd279098080, - 64'd311396925440, 64'd19731441664, 64'd2216447744, - 64'd281278016, - 64'd301096992768, 64'd21449154560, 64'd2029865600, - 64'd282285504, - 64'd289967308800, 64'd23049652224, 64'd1839584256, - 64'd282146208, - 64'd278067412992, 64'd24529580032, 64'd1646428544, - 64'd280889568, - 64'd265458302976, 64'd25886117888, 64'd1451213696, - 64'd278548480, - 64'd252202254336, 64'd27116988416, 64'd1254742784, - 64'd275159200, - 64'd238362558464, 64'd28220442624, 64'd1057803904, - 64'd270761088, - 64'd224003260416, 64'd29195257856, 64'd861167552, - 64'd265396368, - 64'd209188864000, 64'd30040733696, 64'd665584192, - 64'd259109872, - 64'd193984118784, 64'd30756673536, 64'd471781696, - 64'd251948880, - 64'd178453741568, 64'd31343376384, 64'd280463328, - 64'd243962800, - 64'd162662154240, 64'd31801628672, 64'd92305616, - 64'd235202960, - 64'd146673319936, 64'd32132683776, - 64'd92043536, - 64'd225722400, - 64'd130550407168, 64'd32338247680, - 64'd271966656, - 64'd215575552, - 64'd114355642368, 64'd32420460544, - 64'd446878272, - 64'd204818064, - 64'd98150088704, 64'd32381878272, - 64'd616226368, - 64'd193506512, - 64'd81993424896, 64'd32225458176, - 64'd779493568, - 64'd181698208, - 64'd65943736320, 64'd31954526208, - 64'd936198400, - 64'd169450944, - 64'd50057383936, 64'd31572770816, - 64'd1085896192, - 64'd156822736, - 64'd34388787200, 64'd31084206080, - 64'd1228179712, - 64'd143871632, - 64'd18990278656, 64'd30493153280, - 64'd1362680064, - 64'd130655464, - 64'd3911964416, 64'd29804226560, - 64'd1489066880, - 64'd117231656, 64'd10798425088, 64'd29022289920, - 64'd1607048832, - 64'd103657016, 64'd25095653376, 64'd28152449024, - 64'd1716373632, - 64'd89987512, 64'd38937088000, 64'd27200020480, - 64'd1816828288, - 64'd76278104, 64'd52282806272, 64'd26170503168, - 64'd1908238464, - 64'd62582548, 64'd65095667712, 64'd25069555712, - 64'd1990468736, - 64'd48953224, 64'd77341401088, 64'd23902976000, - 64'd2063421824, - 64'd35440968, 64'd88988663808, 64'd22676664320, - 64'd2127038208, - 64'd22094926, 64'd100009091072, 64'd21396609024, - 64'd2181295360, - 64'd8962404, 64'd110377304064, 64'd20068861952, - 64'd2226206464, 64'd3911272, 64'd120070995968, 64'd18699503616, - 64'd2261820928, 64'd16482871, 64'd129070874624, 64'd17294628864, - 64'd2288220928, 64'd28711376, 64'd137360703488, 64'd15860324352, - 64'd2305523200, 64'd40558076, 64'd144927277056, 64'd14402635776, - 64'd2313874944, 64'd51986672, 64'd151760420864, 64'd12927555584, - 64'd2313454848, 64'd62963336, 64'd157852909568, 64'd11441000448, - 64'd2304470016, 64'd73456800, 64'd163200466944, 64'd9948783616, - 64'd2287154944, 64'd83438384, 64'd167801683968, 64'd8456606208, - 64'd2261771008, 64'd92882072, 64'd171657986048, 64'd6970028032, - 64'd2228602624, 64'd101764536, 64'd174773534720, 64'd5494456832, - 64'd2187958272, 64'd110065144, 64'd177155129344, 64'd4035129088, - 64'd2140166272, 64'd117765976, 64'd178812190720, 64'd2597094656, - 64'd2085574912, 64'd124851848, 64'd179756580864, 64'd1185201920, - 64'd2024549248, 64'd131310280, 64'd180002521088, - 64'd195915488, - 64'd1957470464, 64'd137131472, 64'd179566510080, - 64'd1541850496, - 64'd1884733440, 64'd142308320, 64'd178467209216, - 64'd2848434688, - 64'd1806744704, 64'd146836288, 64'd176725278720, - 64'd4111747072, - 64'd1723921280, 64'd150713488, 64'd174363279360, - 64'd5328124416, - 64'd1636688256, 64'd153940496, 64'd171405541376, - 64'd6494167040, - 64'd1545477248, 64'd156520384, 64'd167878017024, - 64'd7606746624, - 64'd1450724736, 64'd158458592, 64'd163808182272, - 64'd8663012352, - 64'd1352869760, 64'd159762848, 64'd159224823808, - 64'd9660390400, - 64'd1252353024, 64'd160443152, 64'd154157973504, - 64'd10596594688, - 64'd1149614208, 64'd160511616, 64'd148638744576, - 64'd11469620224, - 64'd1045091264, 64'd159982336, 64'd142699167744, - 64'd12277748736, - 64'd939218176, 64'd158871408, 64'd136372060160, - 64'd13019549696, - 64'd832423680, 64'd157196688, 64'd129690869760, - 64'd13693872128, - 64'd725129664, 64'd154977808, 64'd122689576960, - 64'd14299848704, - 64'd617749760, 64'd152235920, 64'd115402514432, - 64'd14836889600, - 64'd510688032, 64'd148993680, 64'd107864236032, - 64'd15304677376, - 64'd404337664, 64'd145275136, 64'd100109393920, - 64'd15703163904, - 64'd299079680, 64'd141105488, 64'd92172591104, - 64'd16032561152, - 64'd195281808, 64'd136511104, 64'd84088274944, - 64'd16293335040, - 64'd93297480, 64'd131519288, 64'd75890581504, - 64'd16486198272, 64'd6535211, 64'd126158216, 64'd67613241344, - 64'd16612102144, 64'd103894424, 64'd120456760, 64'd59289448448, - 64'd16672225280, 64'd198475360, 64'd114444408, 64'd50951753728, - 64'd16667965440, 64'd289991040, 64'd108151112, 64'd42631954432, - 64'd16600927232, 64'd378172928, 64'd101607160, 64'd34360999936, - 64'd16472913920, 64'd462771488, 64'd94843072, 64'd26168883200, - 64'd16285911040, 64'd543556672, 64'd87889448, 64'd18084569088, - 64'd16042079232, 64'd620318464, 64'd80776896, 64'd10135899136, - 64'd15743739904, 64'd692866816, 64'd73535864, 64'd2349513216, - 64'd15393361920, 64'd761032320, 64'd66196568, - 64'd5249213952, - 64'd14993550336, 64'd824666176, 64'd58788864, - 64'd12636242944, - 64'd14547033088, 64'd883640000, 64'd51342156, - 64'd19788924928, - 64'd14056644608, 64'd937846208, 64'd43885276, - 64'd26686052352, - 64'd13525316608, 64'd987197824, 64'd36446412, - 64'd33307910144, - 64'd12956062720, 64'd1031628032, 64'd29053004, - 64'd39636299776, - 64'd12351965184, 64'd1071090304, 64'd21731660, - 64'd45654581248, - 64'd11716163584, 64'd1105557888, 64'd14508074, - 64'd51347697664, - 64'd11051837440, 64'd1135023360, 64'd7406957, - 64'd56702189568, - 64'd10362195968, 64'd1159498496, 64'd451962, - 64'd61706203136, - 64'd9650468864, 64'd1179013376, - 64'd6334379, - 64'd66349502464, - 64'd8919883776, 64'd1193616128, - 64'd12930710, - 64'd70623469568, - 64'd8173664768, 64'd1203372032, - 64'd19316906, - 64'd74521083904, - 64'd7415013888, 64'd1208363136, - 64'd25474120, - 64'd78036934656, - 64'd6647101952, 64'd1208687616, - 64'd31384818, - 64'd81167155200, - 64'd5873056768, 64'd1204458240, - 64'd37032824, - 64'd83909468160, - 64'd5095951872, 64'd1195802752, - 64'd42403336, - 64'd86263095296, - 64'd4318798848, 64'd1182862208, - 64'd47482952, - 64'd88228741120, - 64'd3544532992, 64'd1165790336, - 64'd52259696, - 64'd89808576512, - 64'd2776008448, 64'd1144752512, - 64'd56723012, - 64'd91006156800, - 64'd2015987200, 64'd1119925504, - 64'd60863792, - 64'd91826413568, - 64'd1267131008, 64'd1091495424, - 64'd64674348, - 64'd92275572736, - 64'd531994752, 64'd1059657728, - 64'd68148424, - 64'd92361097216, 64'd186981552, 64'd1024616000, - 64'd71281200, - 64'd92091662336, 64'd887478528, 64'd986580736, - 64'd74069224, - 64'd91477065728, 64'd1567303552, 64'd945768640, - 64'd76510448, - 64'd90528145408, 64'd2224395776, 64'd902401664, - 64'd78604176, - 64'd89256771584, 64'd2856830720, 64'd856705792, - 64'd80351032, - 64'd87675723776, 64'd3462824192, 64'd808910336, - 64'd81752936, - 64'd85798625280, 64'd4040735232, 64'd759246976, - 64'd82813040, - 64'd83639910400, 64'd4589070336, 64'd707948672, - 64'd83535736, - 64'd81214709760, 64'd5106482176, 64'd655248832, - 64'd83926560, - 64'd78538784768, 64'd5591775744, 64'd601380672, - 64'd83992160, - 64'd75628462080, 64'd6043904512, 64'd546575744, - 64'd83740256, - 64'd72500551680, 64'd6461974528, 64'd491063776, - 64'd83179568, - 64'd69172289536, 64'd6845240832, 64'd435071360, - 64'd82319768, - 64'd65661214720, 64'd7193108992, 64'd378821440, - 64'd81171424, - 64'd61985153024, 64'd7505132544, 64'd322532448, - 64'd79745920, - 64'd58162106368, 64'd7781011968, 64'd266417632, - 64'd78055424, - 64'd54210191360, 64'd8020591616, 64'd210684352, - 64'd76112784, - 64'd50147569664, 64'd8223855104, 64'd155533488, - 64'd73931496, - 64'd45992374272, 64'd8390925824, 64'd101158768, - 64'd71525640, - 64'd41762639872, 64'd8522059264, 64'd47746272, - 64'd68909760, - 64'd37476241408, 64'd8617641984, - 64'd4526102, - 64'd66098868, - 64'd33150840832, 64'd8678182912, - 64'd55489112, - 64'd63108336, - 64'd28803799040, 64'd8704313344, - 64'd104982600, - 64'd59953832, - 64'd24452141056, 64'd8696778752, - 64'd152855856, - 64'd56651264, - 64'd20112492544, 64'd8656432128, - 64'd198967984, - 64'd53216712, - 64'd15801023488, 64'd8584230912, - 64'd243188192, - 64'd49666348, - 64'd11533401088, 64'd8481228800, - 64'd285396000, - 64'd46016400, - 64'd7324742656, 64'd8348569600, - 64'd325481472, - 64'd42283064, - 64'd3189574144, 64'd8187483136, - 64'd363345376, - 64'd38482464, 64'd858214400, 64'd7999273472, - 64'd398899296, - 64'd34630572};
	localparam logic signed[63:0] hb[0:1199] = {64'd5880330321920, 64'd9331200000, - 64'd12121982976, - 64'd37615036, 64'd5871003762688, 64'd27963885568, - 64'd12043516928, - 64'd112520208, 64'd5852380528640, 64'd46507737088, - 64'd11887098880, - 64'd186471232, 64'd5824520388608, 64'd64904146944, - 64'd11653682176, - 64'd258876112, 64'd5787510374400, 64'd83095248896, - 64'd11344629760, - 64'd329181408, 64'd5741467926528, 64'd101024178176, - 64'd10961692672, - 64'd396872800, 64'd5686538797056, 64'd118635307008, - 64'd10506989568, - 64'd461475424, 64'd5622894428160, 64'd135874502656, - 64'd9982984192, - 64'd522554208, 64'd5550734573568, 64'd152689360896, - 64'd9392459776, - 64'd579713856, 64'd5470283628544, 64'd169029353472, - 64'd8738495488, - 64'd632598976, 64'd5381791678464, 64'd184846123008, - 64'd8024443392, - 64'd680893760, 64'd5285531877376, 64'd200093564928, - 64'd7253902336, - 64'd724321536, 64'd5181799923712, 64'd214728081408, - 64'd6430694400, - 64'd762644672, 64'd5070912487424, 64'd228708646912, - 64'd5558839296, - 64'd795663808, 64'd4953206685696, 64'd241997037568, - 64'd4642529792, - 64'd823217088, 64'd4829036412928, 64'd254557880320, - 64'd3686106112, - 64'd845179392, 64'd4698774962176, 64'd266358784000, - 64'd2694032896, - 64'd861461696, 64'd4562809257984, 64'd277370437632, - 64'd1670873728, - 64'd872009664, 64'd4421540380672, 64'd287566626816, - 64'd621268032, - 64'd876802624, 64'd4275381993472, 64'd296924446720, 64'd450092960, - 64'd875852672, 64'd4124758769664, 64'd305424171008, 64'd1538488960, - 64'd869203008, 64'd3970103508992, 64'd313049317376, 64'd2639193088, - 64'd856926848, 64'd3811857137664, 64'd319786811392, 64'd3747492864, - 64'd839125696, 64'd3650466086912, 64'd325626822656, 64'd4858712576, - 64'd815928384, 64'd3486380982272, 64'd330562732032, 64'd5968231424, - 64'd787488832, 64'd3320054546432, 64'd334591328256, 64'd7071505408, - 64'd753985088, 64'd3151940812800, 64'd337712480256, 64'd8164083712, - 64'd715617280, 64'd2982492766208, 64'd339929333760, 64'd9241626624, - 64'd672606272, 64'd2812161032192, 64'd341248049152, 64'd10299923456, - 64'd625191680, 64'd2641392828416, 64'd341677899776, 64'd11334905856, - 64'd573630336, 64'd2470629343232, 64'd341231042560, 64'd12342664192, - 64'd518194528, 64'd2300305211392, 64'd339922550784, 64'd13319460864, - 64'd459170304, 64'd2130847334400, 64'd337770184704, 64'd14261741568, - 64'd396855712, 64'd1962672390144, 64'd334794358784, 64'd15166146560, - 64'd331559072, 64'd1796186439680, 64'd331017977856, 64'd16029522944, - 64'd263597264, 64'd1631783616512, 64'd326466371584, 64'd16848930816, - 64'd193294128, 64'd1469844684800, 64'd321167097856, 64'd17621653504, - 64'd120978672, 64'd1310736252928, 64'd315149746176, 64'd18345203712, - 64'd46983556, 64'd1154809462784, 64'd308446003200, 64'd19017326592, 64'd28356576, 64'd1002399203328, 64'd301089226752, 64'd19636006912, 64'd104706624, 64'd853823324160, 64'd293114478592, 64'd20199477248, 64'd181732544, 64'd709381718016, 64'd284558295040, 64'd20706205696, 64'd259102800, 64'd569355730944, 64'd275458523136, 64'd21154916352, 64'd336489792, 64'd434007375872, 64'd265854238720, 64'd21544572928, 64'd413571200, 64'd303579004928, 64'd255785402368, 64'd21874386944, 64'd490031264, 64'd178292686848, 64'd245292875776, 64'd22143815680, 64'd565561984, 64'd58349928448, 64'd234418176000, 64'd22352556032, 64'd639864384, - 64'd56068689920, 64'd223203344384, 64'd22500540416, 64'd712649344, - 64'd164803657728, 64'd211690684416, 64'd22587938816, 64'd783638912, - 64'd267716722688, 64'd199922761728, 64'd22615146496, 64'd852567168, - 64'd364690866176, 64'd187942109184, 64'd22582779904, 64'd919180992, - 64'd455630323712, 64'd175791144960, 64'd22491672576, 64'd983240768, - 64'd540460515328, 64'd163512008704, 64'd22342860800, 64'd1044521472, - 64'd619127832576, 64'd151146397696, 64'd22137585664, 64'd1102812928, - 64'd691599245312, 64'd138735403008, 64'd21877274624, 64'd1157920384, - 64'd757862301696, 64'd126319476736, 64'd21563535360, 64'd1209665408, - 64'd817924407296, 64'd113938153472, 64'd21198149632, 64'd1257885696, - 64'd871812562944, 64'd101630058496, 64'd20783056896, 64'd1302435840, - 64'd919572840448, 64'd89432686592, 64'd20320348160, 64'd1343187328, - 64'd961269661696, 64'd77382361088, 64'd19812251648, 64'd1380028928, - 64'd996985405440, 64'd65514090496, 64'd19261124608, 64'd1412866432, - 64'd1026819620864, 64'd53861486592, 64'd18669438976, 64'd1441623168, - 64'd1050888110080, 64'd42456657920, 64'd18039771136, 64'd1466239488, - 64'd1069322600448, 64'd31330148352, 64'd17374785536, 64'd1486672896, - 64'd1082269433856, 64'd20510838784, 64'd16677234688, 64'd1502897792, - 64'd1089889107968, 64'd10025896960, 64'd15949931520, 64'd1514905216, - 64'd1092355227648, - 64'd99294480, 64'd15195747328, 64'd1522702848, - 64'd1089853652992, - 64'd9841181696, 64'd14417598464, 64'd1526313984, - 64'd1082581450752, - 64'd19178088448, 64'd13618429952, 64'd1525777664, - 64'd1070746304512, - 64'd28090251264, 64'd12801209344, 64'd1521148160, - 64'd1054564941824, - 64'd36559847424, 64'd11968911360, 64'd1512493952, - 64'd1034262806528, - 64'd44571013120, 64'd11124508672, 64'd1499897856, - 64'd1010072616960, - 64'd52109860864, 64'd10270958592, 64'd1483456128, - 64'd982233645056, - 64'd59164479488, 64'd9411194880, 64'd1463277440, - 64'd950990536704, - 64'd65724940288, 64'd8548114432, 64'd1439482880, - 64'd916592394240, - 64'd71783268352, 64'd7684571136, 64'd1412204416, - 64'd879291924480, - 64'd77333463040, 64'd6823361024, 64'd1381585280, - 64'd839344324608, - 64'd82371428352, 64'd5967217664, 64'd1347777792, - 64'd797006233600, - 64'd86894968832, 64'd5118800896, 64'd1310943872, - 64'd752535142400, - 64'd90903748608, 64'd4280687872, 64'd1271253504, - 64'd706188083200, - 64'd94399275008, 64'd3455368448, 64'd1228883712, - 64'd658220908544, - 64'd97384783872, 64'd2645234176, 64'd1184018688, - 64'd608887504896, - 64'd99865255936, 64'd1852573824, 64'd1136848000, - 64'd558438744064, - 64'd101847326720, 64'd1079566336, 64'd1087566080, - 64'd507121893376, - 64'd103339220992, 64'd328275104, 64'd1036371520, - 64'd455179632640, - 64'd104350679040, - 64'd399356832, 64'd983466112, - 64'd402849431552, - 64'd104892923904, - 64'd1101511680, 64'd929053952, - 64'd350362861568, - 64'd104978538496, - 64'd1776500480, 64'd873340736, - 64'd297944743936, - 64'd104621391872, - 64'd2422767104, 64'd816532992, - 64'd245812789248, - 64'd103836614656, - 64'd3038890496, 64'd758836928, - 64'd194176761856, - 64'd102640427008, - 64'd3623587072, 64'd700458176, - 64'd143238103040, - 64'd101050114048, - 64'd4175712512, 64'd641600704, - 64'd93189341184, - 64'd99083935744, - 64'd4694262784, 64'd582466112, - 64'd44213682176, - 64'd96760987648, - 64'd5178375168, 64'd523253056, 64'd3515442688, - 64'd94101176320, - 64'd5627326976, 64'd464156384, 64'd49834721280, - 64'd91125080064, - 64'd6040537088, 64'd405366656, 64'd94591270912, - 64'd87853858816, - 64'd6417562624, 64'd347069472, 64'd137642950656, - 64'd84309204992, - 64'd6758099456, 64'd289444800, 64'd178858524672, - 64'd80513187840, - 64'd7061979136, 64'd232666592, 64'd218117931008, - 64'd76488237056, - 64'd7329165824, 64'd176902112, 64'd255312314368, - 64'd72256970752, - 64'd7559755264, 64'd122311512, 64'd290344239104, - 64'd67842166784, - 64'd7753970176, 64'd69047432, 64'd323127640064, - 64'd63266664448, - 64'd7912156160, 64'd17254548, 64'd353587888128, - 64'd58553266176, - 64'd8034778112, - 64'd32930780, 64'd381661642752, - 64'd53724651520, - 64'd8122417152, - 64'd81380816, 64'd407297032192, - 64'd48803319808, - 64'd8175762432, - 64'd127976752, 64'd430453161984, - 64'd43811487744, - 64'd8195609600, - 64'd172608928, 64'd451100344320, - 64'd38771027968, - 64'd8182854144, - 64'd215177056, 64'd469219639296, - 64'd33703397376, - 64'd8138483712, - 64'd255590368, 64'd484802691072, - 64'd28629559296, - 64'd8063577088, - 64'd293767776, 64'd497851531264, - 64'd23569926144, - 64'd7959292416, - 64'd329637856, 64'd508378251264, - 64'd18544300032, - 64'd7826866176, - 64'd363139040, 64'd516404641792, - 64'd13571805184, - 64'd7667602432, - 64'd394219488, 64'd521961930752, - 64'd8670844928, - 64'd7482871296, - 64'd422837184, 64'd525090324480, - 64'd3859045632, - 64'd7274096640, - 64'd448959712, 64'd525838614528, 64'd846788480, - 64'd7042754560, - 64'd472564352, 64'd524263817216, 64'd5430713856, - 64'd6790364160, - 64'd493637728, 64'd520430714880, 64'd9877687296, - 64'd6518481408, - 64'd512175872, 64'd514411298816, 64'd14173598720, - 64'd6228693504, - 64'd528183840, 64'd506284474368, 64'd18305296384, - 64'd5922609664, - 64'd541675520, 64'd496135405568, 64'd22260619264, - 64'd5601858560, - 64'd552673600, 64'd484055089152, 64'd26028408832, - 64'd5268078080, - 64'd561208832, 64'd470139928576, 64'd29598525440, - 64'd4922912768, - 64'd567320192, 64'd454491045888, 64'd32961867776, - 64'd4568003584, - 64'd571054272, 64'd437213855744, 64'd36110372864, - 64'd4204985344, - 64'd572465024, 64'd418417639424, 64'd39037022208, - 64'd3835479296, - 64'd571613376, 64'd398214823936, 64'd41735839744, - 64'd3461087744, - 64'd568566912, 64'd376720621568, 64'd44201889792, - 64'd3083388160, - 64'd563399296, 64'd354052407296, 64'd46431268864, - 64'd2703929344, - 64'd556190080, 64'd330329292800, 64'd48421093376, - 64'd2324225024, - 64'd547024064, 64'd305671569408, 64'd50169475072, - 64'd1945749504, - 64'd535990976, 64'd280200216576, 64'd51675516928, - 64'd1569933696, - 64'd523185088, 64'd254036443136, 64'd52939288576, - 64'd1198160256, - 64'd508704608, 64'd227301163008, 64'd53961793536, - 64'd831760256, - 64'd492651296, 64'd200114569216, 64'd54744944640, - 64'd472009056, - 64'd475130048, 64'd172595675136, 64'd55291535360, - 64'd120123344, - 64'd456248384, 64'd144861888512, 64'd55605202944, 64'd222742160, - 64'd436116000, 64'd117028585472, 64'd55690399744, 64'd555497280, - 64'd414844320, 64'd89208733696, 64'd55552348160, 64'd877118976, - 64'd392546016, 64'd61512495104, 64'd55196999680, 64'd1186653184, - 64'd369334656, 64'd34046879744, 64'd54631010304, 64'd1483216768, - 64'd345324096, 64'd6915413504, 64'd53861675008, 64'd1765999360, - 64'd320628256, - 64'd19782180864, 64'd52896890880, 64'd2034263808, - 64'd295360544, - 64'd45950271488, 64'd51745124352, 64'd2287347712, - 64'd269633472, - 64'd71497596928, 64'd50415345664, 64'd2524663808, - 64'd243558400, - 64'd96337477632, 64'd48916996096, 64'd2745700096, - 64'd217244960, - 64'd120388091904, 64'd47259926528, 64'd2950020096, - 64'd190800800, - 64'd143572615168, 64'd45454368768, 64'd3137262336, - 64'd164331248, - 64'd165819432960, 64'd43510865920, 64'd3307140096, - 64'd137938944, - 64'd187062255616, 64'd41440239616, 64'd3459440128, - 64'd111723488, - 64'd207240282112, 64'd39253532672, 64'd3594022400, - 64'd85781248, - 64'd226298265600, 64'd36961959936, 64'd3710817792, - 64'd60205020, - 64'd244186611712, 64'd34576879616, 64'd3809826816, - 64'd35083764, - 64'd260861427712, 64'd32109721600, 64'd3891118848, - 64'd10502396, - 64'd276284538880, 64'd29571948544, 64'd3954828288, 64'd13458433, - 64'd290423472128, 64'd26975027200, 64'd4001154304, 64'd36722532, - 64'd303251554304, 64'd24330364928, 64'd4030357248, 64'd59218340, - 64'd314747748352, 64'd21649278976, 64'd4042756096, 64'd80879072, - 64'd324896587776, 64'd18942945280, 64'd4038726400, 64'd101642872, - 64'd333688274944, 64'd16222372864, 64'd4018696960, 64'd121452864, - 64'd341118353408, 64'd13498356736, 64'd3983147776, 64'd140257312, - 64'd347187773440, 64'd10781442048, 64'd3932604928, 64'd158009632, - 64'd351902662656, 64'd8081892864, 64'd3867639552, 64'd174668432, - 64'd355274194944, 64'd5409659904, 64'd3788863488, 64'd190197584, - 64'd357318459392, 64'd2774347008, 64'd3696925696, 64'd204566176, - 64'd358056230912, 64'd185187008, 64'd3592510208, 64'd217748528, - 64'd357512806400, - 64'd2348986880, 64'd3476330752, 64'd229724128, - 64'd355717775360, - 64'd4819764224, 64'd3349128448, 64'd240477616, - 64'd352704888832, - 64'd7219179520, 64'd3211668736, 64'd249998672, - 64'd348511731712, - 64'd9539730432, 64'd3064736512, 64'd258281952, - 64'd343179460608, - 64'd11774398464, 64'd2909133824, 64'd265326992, - 64'd336752738304, - 64'd13916656640, 64'd2745675776, 64'd271138016, - 64'd329279209472, - 64'd15960493056, 64'd2575187456, 64'd275723936, - 64'd320809533440, - 64'd17900410880, 64'd2398499840, 64'd279098080, - 64'd311396925440, - 64'd19731441664, 64'd2216447744, 64'd281278016, - 64'd301096992768, - 64'd21449154560, 64'd2029865600, 64'd282285504, - 64'd289967308800, - 64'd23049652224, 64'd1839584256, 64'd282146208, - 64'd278067412992, - 64'd24529580032, 64'd1646428544, 64'd280889568, - 64'd265458302976, - 64'd25886117888, 64'd1451213696, 64'd278548480, - 64'd252202254336, - 64'd27116988416, 64'd1254742784, 64'd275159200, - 64'd238362558464, - 64'd28220442624, 64'd1057803904, 64'd270761088, - 64'd224003260416, - 64'd29195257856, 64'd861167552, 64'd265396368, - 64'd209188864000, - 64'd30040733696, 64'd665584192, 64'd259109872, - 64'd193984118784, - 64'd30756673536, 64'd471781696, 64'd251948880, - 64'd178453741568, - 64'd31343376384, 64'd280463328, 64'd243962800, - 64'd162662154240, - 64'd31801628672, 64'd92305616, 64'd235202960, - 64'd146673319936, - 64'd32132683776, - 64'd92043536, 64'd225722400, - 64'd130550407168, - 64'd32338247680, - 64'd271966656, 64'd215575552, - 64'd114355642368, - 64'd32420460544, - 64'd446878272, 64'd204818064, - 64'd98150088704, - 64'd32381878272, - 64'd616226368, 64'd193506512, - 64'd81993424896, - 64'd32225458176, - 64'd779493568, 64'd181698208, - 64'd65943736320, - 64'd31954526208, - 64'd936198400, 64'd169450944, - 64'd50057383936, - 64'd31572770816, - 64'd1085896192, 64'd156822736, - 64'd34388787200, - 64'd31084206080, - 64'd1228179712, 64'd143871632, - 64'd18990278656, - 64'd30493153280, - 64'd1362680064, 64'd130655464, - 64'd3911964416, - 64'd29804226560, - 64'd1489066880, 64'd117231656, 64'd10798425088, - 64'd29022289920, - 64'd1607048832, 64'd103657016, 64'd25095653376, - 64'd28152449024, - 64'd1716373632, 64'd89987512, 64'd38937088000, - 64'd27200020480, - 64'd1816828288, 64'd76278104, 64'd52282806272, - 64'd26170503168, - 64'd1908238464, 64'd62582548, 64'd65095667712, - 64'd25069555712, - 64'd1990468736, 64'd48953224, 64'd77341401088, - 64'd23902976000, - 64'd2063421824, 64'd35440968, 64'd88988663808, - 64'd22676664320, - 64'd2127038208, 64'd22094926, 64'd100009091072, - 64'd21396609024, - 64'd2181295360, 64'd8962404, 64'd110377304064, - 64'd20068861952, - 64'd2226206464, - 64'd3911272, 64'd120070995968, - 64'd18699503616, - 64'd2261820928, - 64'd16482871, 64'd129070874624, - 64'd17294628864, - 64'd2288220928, - 64'd28711376, 64'd137360703488, - 64'd15860324352, - 64'd2305523200, - 64'd40558076, 64'd144927277056, - 64'd14402635776, - 64'd2313874944, - 64'd51986672, 64'd151760420864, - 64'd12927555584, - 64'd2313454848, - 64'd62963336, 64'd157852909568, - 64'd11441000448, - 64'd2304470016, - 64'd73456800, 64'd163200466944, - 64'd9948783616, - 64'd2287154944, - 64'd83438384, 64'd167801683968, - 64'd8456606208, - 64'd2261771008, - 64'd92882072, 64'd171657986048, - 64'd6970028032, - 64'd2228602624, - 64'd101764536, 64'd174773534720, - 64'd5494456832, - 64'd2187958272, - 64'd110065144, 64'd177155129344, - 64'd4035129088, - 64'd2140166272, - 64'd117765976, 64'd178812190720, - 64'd2597094656, - 64'd2085574912, - 64'd124851848, 64'd179756580864, - 64'd1185201920, - 64'd2024549248, - 64'd131310280, 64'd180002521088, 64'd195915488, - 64'd1957470464, - 64'd137131472, 64'd179566510080, 64'd1541850496, - 64'd1884733440, - 64'd142308320, 64'd178467209216, 64'd2848434688, - 64'd1806744704, - 64'd146836288, 64'd176725278720, 64'd4111747072, - 64'd1723921280, - 64'd150713488, 64'd174363279360, 64'd5328124416, - 64'd1636688256, - 64'd153940496, 64'd171405541376, 64'd6494167040, - 64'd1545477248, - 64'd156520384, 64'd167878017024, 64'd7606746624, - 64'd1450724736, - 64'd158458592, 64'd163808182272, 64'd8663012352, - 64'd1352869760, - 64'd159762848, 64'd159224823808, 64'd9660390400, - 64'd1252353024, - 64'd160443152, 64'd154157973504, 64'd10596594688, - 64'd1149614208, - 64'd160511616, 64'd148638744576, 64'd11469620224, - 64'd1045091264, - 64'd159982336, 64'd142699167744, 64'd12277748736, - 64'd939218176, - 64'd158871408, 64'd136372060160, 64'd13019549696, - 64'd832423680, - 64'd157196688, 64'd129690869760, 64'd13693872128, - 64'd725129664, - 64'd154977808, 64'd122689576960, 64'd14299848704, - 64'd617749760, - 64'd152235920, 64'd115402514432, 64'd14836889600, - 64'd510688032, - 64'd148993680, 64'd107864236032, 64'd15304677376, - 64'd404337664, - 64'd145275136, 64'd100109393920, 64'd15703163904, - 64'd299079680, - 64'd141105488, 64'd92172591104, 64'd16032561152, - 64'd195281808, - 64'd136511104, 64'd84088274944, 64'd16293335040, - 64'd93297480, - 64'd131519288, 64'd75890581504, 64'd16486198272, 64'd6535211, - 64'd126158216, 64'd67613241344, 64'd16612102144, 64'd103894424, - 64'd120456760, 64'd59289448448, 64'd16672225280, 64'd198475360, - 64'd114444408, 64'd50951753728, 64'd16667965440, 64'd289991040, - 64'd108151112, 64'd42631954432, 64'd16600927232, 64'd378172928, - 64'd101607160, 64'd34360999936, 64'd16472913920, 64'd462771488, - 64'd94843072, 64'd26168883200, 64'd16285911040, 64'd543556672, - 64'd87889448, 64'd18084569088, 64'd16042079232, 64'd620318464, - 64'd80776896, 64'd10135899136, 64'd15743739904, 64'd692866816, - 64'd73535864, 64'd2349513216, 64'd15393361920, 64'd761032320, - 64'd66196568, - 64'd5249213952, 64'd14993550336, 64'd824666176, - 64'd58788864, - 64'd12636242944, 64'd14547033088, 64'd883640000, - 64'd51342156, - 64'd19788924928, 64'd14056644608, 64'd937846208, - 64'd43885276, - 64'd26686052352, 64'd13525316608, 64'd987197824, - 64'd36446412, - 64'd33307910144, 64'd12956062720, 64'd1031628032, - 64'd29053004, - 64'd39636299776, 64'd12351965184, 64'd1071090304, - 64'd21731660, - 64'd45654581248, 64'd11716163584, 64'd1105557888, - 64'd14508074, - 64'd51347697664, 64'd11051837440, 64'd1135023360, - 64'd7406957, - 64'd56702189568, 64'd10362195968, 64'd1159498496, - 64'd451962, - 64'd61706203136, 64'd9650468864, 64'd1179013376, 64'd6334379, - 64'd66349502464, 64'd8919883776, 64'd1193616128, 64'd12930710, - 64'd70623469568, 64'd8173664768, 64'd1203372032, 64'd19316906, - 64'd74521083904, 64'd7415013888, 64'd1208363136, 64'd25474120, - 64'd78036934656, 64'd6647101952, 64'd1208687616, 64'd31384818, - 64'd81167155200, 64'd5873056768, 64'd1204458240, 64'd37032824, - 64'd83909468160, 64'd5095951872, 64'd1195802752, 64'd42403336, - 64'd86263095296, 64'd4318798848, 64'd1182862208, 64'd47482952, - 64'd88228741120, 64'd3544532992, 64'd1165790336, 64'd52259696, - 64'd89808576512, 64'd2776008448, 64'd1144752512, 64'd56723012, - 64'd91006156800, 64'd2015987200, 64'd1119925504, 64'd60863792, - 64'd91826413568, 64'd1267131008, 64'd1091495424, 64'd64674348, - 64'd92275572736, 64'd531994752, 64'd1059657728, 64'd68148424, - 64'd92361097216, - 64'd186981552, 64'd1024616000, 64'd71281200, - 64'd92091662336, - 64'd887478528, 64'd986580736, 64'd74069224, - 64'd91477065728, - 64'd1567303552, 64'd945768640, 64'd76510448, - 64'd90528145408, - 64'd2224395776, 64'd902401664, 64'd78604176, - 64'd89256771584, - 64'd2856830720, 64'd856705792, 64'd80351032, - 64'd87675723776, - 64'd3462824192, 64'd808910336, 64'd81752936, - 64'd85798625280, - 64'd4040735232, 64'd759246976, 64'd82813040, - 64'd83639910400, - 64'd4589070336, 64'd707948672, 64'd83535736, - 64'd81214709760, - 64'd5106482176, 64'd655248832, 64'd83926560, - 64'd78538784768, - 64'd5591775744, 64'd601380672, 64'd83992160, - 64'd75628462080, - 64'd6043904512, 64'd546575744, 64'd83740256, - 64'd72500551680, - 64'd6461974528, 64'd491063776, 64'd83179568, - 64'd69172289536, - 64'd6845240832, 64'd435071360, 64'd82319768, - 64'd65661214720, - 64'd7193108992, 64'd378821440, 64'd81171424, - 64'd61985153024, - 64'd7505132544, 64'd322532448, 64'd79745920, - 64'd58162106368, - 64'd7781011968, 64'd266417632, 64'd78055424, - 64'd54210191360, - 64'd8020591616, 64'd210684352, 64'd76112784, - 64'd50147569664, - 64'd8223855104, 64'd155533488, 64'd73931496, - 64'd45992374272, - 64'd8390925824, 64'd101158768, 64'd71525640, - 64'd41762639872, - 64'd8522059264, 64'd47746272, 64'd68909760, - 64'd37476241408, - 64'd8617641984, - 64'd4526102, 64'd66098868, - 64'd33150840832, - 64'd8678182912, - 64'd55489112, 64'd63108336, - 64'd28803799040, - 64'd8704313344, - 64'd104982600, 64'd59953832, - 64'd24452141056, - 64'd8696778752, - 64'd152855856, 64'd56651264, - 64'd20112492544, - 64'd8656432128, - 64'd198967984, 64'd53216712, - 64'd15801023488, - 64'd8584230912, - 64'd243188192, 64'd49666348, - 64'd11533401088, - 64'd8481228800, - 64'd285396000, 64'd46016400, - 64'd7324742656, - 64'd8348569600, - 64'd325481472, 64'd42283064, - 64'd3189574144, - 64'd8187483136, - 64'd363345376, 64'd38482464, 64'd858214400, - 64'd7999273472, - 64'd398899296, 64'd34630572};
endpackage
`endif
