`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam real Lfr[0:2] = {0.970789348297097, 0.9498022845398874, 0.9707893482970972};
	localparam real Lfi[0:2] = {0.0813884092055478, -1.7722241656505967e-15, -0.08138840920554608};
	localparam real Lbr[0:2] = {0.9707893482970993, 0.9498022845398779, 0.9707893482971011};
	localparam real Lbi[0:2] = {0.08138840920555224, -3.791305919383092e-15, -0.08138840920554852};
	localparam real Wfr[0:2] = {0.0006240970025894416, -0.0009360490045281465, 0.0006240970025893649};
	localparam real Wfi[0:2] = {-0.0010474400734392735, -1.015051476217961e-18, 0.0010474400734392512};
	localparam real Wbr[0:2] = {-0.0006248243462250154, 0.0009379784791755657, -0.0006248243462248402};
	localparam real Wbi[0:2] = {0.001048491217384701, -5.484447390469192e-18, -0.0010484912173847204};
	localparam real Ffr[0:2][0:59] = '{
		'{8.005326134896476, -0.805739580014779, -0.08456475319940855, 7.54404899082117, -0.8816207661123752, -0.0685024663388227, 7.049861750830094, -0.9470440893890363, -0.052746240195884725, 6.528136189506291, -1.0020531227482206, -0.037398297409506065, 5.98417633518283, -1.0467670904546773, -0.02255260012017933, 5.423182261207181, -1.081376122674106, -0.00829456820611383, 4.850216499128535, -1.106136221578197, 0.005299124253100321, 4.270173191376808, -1.1213639913491789, 0.018160676748610313, 3.6877500745284704, -1.1274311835172925, 0.030231217254536265, 3.107423358448414, -1.1247591078252037, 0.04146078758149849, 2.5334255416175364, -1.1138129572617903, 0.05180826282454957, 1.9697261789472977, -1.0950960940714782, 0.06124120886531876, 1.4200155954753553, -1.0691443414526134, 0.06973568214963716, 0.8876915176455833, -1.0365203233379325, 0.07727597617848928, 0.37584857350151757, -0.9978078921309967, 0.08385431932249836, -0.11272940584999613, -0.9536066815834512, 0.08947052869925957, -0.5755743686482571, -0.9045268191678969, 0.09413162493992956, -1.0105364098764005, -0.8511838293584013, 0.09785141271804816, -1.4157836391645588, -0.7941937562029349, 0.1006500319213267, -1.7897996775204168, -0.7341685304862913, 0.10255348431800555},
		'{-15.714065250214375, 1.4604890833954896, -0.312393945388571, -14.92525507406247, 1.387175867954602, -0.29671248300649355, -14.17604136668508, 1.317542808441882, -0.28181819421107007, -13.464436475809435, 1.2514051694371988, -0.26767156468658004, -12.788552524765992, 1.1885874888164762, -0.25423506364567994, -12.146596403981084, 1.128923112253417, -0.24147304426081048, -11.536865013885215, 1.0722537510881753, -0.22935164909371916, -10.957740746616475, 1.0184290623900125, -0.217838720272205, -10.40768719453214, 0.9673062500998494, -0.20690371417578582, -9.885245074143157, 0.9187496861945487, -0.19651762040394924, -9.38902835465784, 0.872630550867887, -0.1866528848120134, -8.917720580863795, 0.8288264907736194, -0.17728333641041075, -8.470071380592804, 0.7872212944239616, -0.16838411793346153, -8.044893147502963, 0.7477045838823259, -0.15993161989343554, -7.641057890377601, 0.7101715219323791, -0.15190341794495002, -7.257494240582176, 0.6745225339465424, -0.14427821339353084, -6.893184609740026, 0.6406630437160596, -0.13703577669050895, -6.547162490086269, 0.6085032225417911, -0.13015689376434325, -6.218509890337796, 0.5779577509200768, -0.12362331504598865, -5.906354900276723, 0.548945592191424, -0.11741770705307424},
		'{8.005326134896897, -0.8057395800148376, -0.08456475319940303, 7.544048990821559, -0.8816207661124327, -0.06850246633881739, 7.049861750830452, -0.9470440893890928, -0.05274624019587969, 6.528136189506619, -1.0020531227482758, -0.03739829740950132, 5.98417633518313, -1.0467670904547313, -0.02255260012017491, 5.423182261207452, -1.081376122674159, -0.00829456820610975, 4.850216499128779, -1.1061362215782484, 0.005299124253104054, 4.270173191377026, -1.121363991349229, 0.018160676748613665, 3.687750074528662, -1.1274311835173414, 0.030231217254539255, 3.107423358448581, -1.1247591078252515, 0.04146078758150112, 2.53342554161768, -1.1138129572618367, 0.05180826282455185, 1.9697261789474168, -1.0950960940715235, 0.06124120886532073, 1.4200155954754536, -1.0691443414526578, 0.0697356821496388, 0.8876915176456588, -1.0365203233379758, 0.07727597617849066, 0.3758485735015724, -0.9978078921310392, 0.0838543193224995, -0.11272940584996172, -0.9536066815834925, 0.08947052869926049, -0.5755743686482424, -0.9045268191679371, 0.0941316249399303, -1.010536409876405, -0.8511838293584407, 0.09785141271804876, -1.4157836391645817, -0.7941937562029732, 0.10065003192132715, -1.7897996775204577, -0.7341685304863286, 0.10255348431800591}};
localparam real Ffi[0:2][0:59] = '{
	'{2.7944562721001764, 1.2215174777721856, -0.16700283788824172, 3.364369142527686, 1.1202582935286247, -0.16900716689505155, 3.8800918736369683, 1.0157811070226088, -0.16964566416955912, 4.340528894359993, 0.9090310670160917, -0.16898313634171125, 4.7450538361615395, 0.8009221675304371, -0.16709081673552498, 5.093490313567917, 0.6923320007527455, -0.1640455053323402, 5.386090319137572, 0.5840970494386741, -0.15992871092399297, 5.6235105159514385, 0.4770085265279428, -0.1548258017587556, 5.8067867120007035, 0.3718087652039268, -0.14882517059829228, 5.937306799956918, 0.26918815834826804, -0.14201741969462645, 6.016782442842376, 0.16978264228686635, -0.13449457076651442, 6.047219781205319, 0.0741717159137622, -0.1263493046089293, 6.030889430680668, -0.017123017269688068, -0.11767423451172085, 5.970296030425143, -0.10363879993806163, -0.10856121719797056, 5.868147593003601, -0.1849721832758584, -0.09910070452298436, 5.7273248950226066, -0.26077902228874444, -0.08938113870497899, 5.550851135311918, -0.33077402791910265, -0.07948839339184693, 5.341862073899888, -0.3947299018930207, -0.06950526240826022, 5.103576850570125, -0.4524760820250693, -0.059510997576896194, 4.839269666578277, -0.5038971272074764, -0.04958089656962079},
	'{3.180953950060241e-13, 3.1578057303335035e-14, -3.1492050425864598e-15, 3.2997657905537974e-13, 2.7404596920776717e-14, -2.4374900447125944e-15, 3.3986340635220914e-13, 2.3570562167052e-14, -1.7892925803769547e-15, 3.479261628681381e-13, 2.0052392589755567e-14, -1.2000291664514298e-15, 3.5432306404265135e-13, 1.6828037809943865e-14, -6.654164284150009e-16, 3.592010375209653e-13, 1.3876865285537767e-14, -1.8145252033034828e-16, 3.626964577240506e-13, 1.1179573529759041e-14, 2.556003460469387e-16, 3.6493583511428417e-13, 8.718110469358826e-15, 6.49232327560273e-16, 3.660364628541067e-13, 6.475596645299664e-15, 1.0027013921946983e-15, 3.6610702339841227e-13, 4.436252975452637e-15, 1.3190478352430413e-15, 3.6524815741368503e-13, 2.5853328148239073e-15, 1.6011079231872636e-15, 3.6355299727760574e-13, 9.090580638826237e-16, 1.8515267162904247e-15, 3.611076672815199e-13, -6.054409102252692e-16, 2.072770117972976e-15, 3.5799175253432915e-13, -1.9701817613787574e-15, 2.2671361962901843e-15, 3.542787384496255e-13, -3.1963832702403417e-15, 2.43676582022628e-15, 3.5003642258782587e-13, -4.29451526526478e-15, 2.5836526510665956e-15, 3.453273005213162e-13, -5.274345544875846e-15, 2.7096525267934986e-15, 3.4020892729281047e-13, -6.144983976088722e-15, 2.816492275267362e-15, 3.3473425594494783e-13, -6.914923934814891e-15, 2.905777989893072e-15, 3.2895195451226463e-13, -7.59208124361236e-15, 2.9790027995284994e-15},
	'{-2.7944562721004997, -1.2215174777722173, 0.16700283788824485, -3.364369142528021, -1.1202582935286525, 0.16900716689505402, -3.880091873637313, -1.0157811070226328, 0.16964566416956103, -4.340528894360347, -0.9090310670161125, 0.16898313634171266, -4.745053836161899, -0.8009221675304548, 0.16709081673552595, -5.093490313568281, -0.69233200075276, 0.16404550533234077, -5.386090319137939, -0.5840970494386861, 0.15992871092399324, -5.623510515951808, -0.4770085265279522, 0.15482580175875557, -5.806786712001074, -0.3718087652039339, 0.1488251705982921, -5.9373067999572875, -0.269188158348273, 0.14201741969462606, -6.016782442842744, -0.16978264228686935, 0.13449457076651394, -6.047219781205685, -0.0741717159137632, 0.12634930460892876, -6.0308894306810314, 0.017123017269688623, 0.11767423451172035, -5.970296030425503, 0.10363879993806407, 0.10856121719797007, -5.8681475930039575, 0.1849721832758625, 0.09910070452298395, -5.727324895022957, 0.2607790222887502, 0.08938113870497866, -5.5508511353122625, 0.3307740279191101, 0.07948839339184671, -5.341862073900226, 0.3947299018930298, 0.06950526240826012, -5.103576850570456, 0.45247608202507994, 0.059510997576896235, -4.8392696665786, 0.5038971272074885, 0.04958089656962098}};
	localparam real Fbr[0:2][0:59] = '{
		'{-7.997160167675694, -0.964793223786971, 0.06746783761726301, -7.53640548355534, -1.0313925870869098, 0.049983942051988944, -7.0427712404028355, -1.0868870463224407, 0.03301699880867022, -6.521623522188401, -1.131427378691316, 0.016667539808804407, -5.978260770750787, -1.1652385878823242, 0.00102635834214259, -5.41787761352952, -1.1886144402552672, -0.013825673700638696, -4.845531310311087, -1.2019117652080653, -0.027817705098744747, -4.2661109364550205, -1.205544574362293, -0.04088892458691212, -3.684309393620068, -1.1999780527700783, -0.05298850408645663, -3.104598313231597, -1.185722473591869, -0.06407547018072308, -2.5312058929776766, -1.1633270856457505, -0.07411850845147332, -1.9680976826376837, -1.1333740209151988, -0.08309570555958481, -1.4189603126635255, -1.0964722665541073, -0.09099423417016106, -0.8871881372648476, -1.0532517431766841, -0.0978099859897066, -0.3758727433959417, -1.0043575282962554, -0.10354715830264838, 0.11220474191119822, -0.9504442607118044, -0.10821779946773599, 0.5745786309059133, -0.8921707584643209, -0.11184131886354351, 1.0091010421643198, -0.8301948797262194, -0.11444396675847845, 1.4139417707035873, -0.7651686526747008, -0.11605828952664926, 1.7875857893398401, -0.69773369706152, -0.11672256553910443},
		'{15.68174053148843, 1.770984996776288, 0.34471540725882666, 14.89455298236931, 1.6820855958239667, 0.327411481330528, 14.146880449854622, 1.5976487417052252, 0.31097617295232105, 13.436739370384457, 1.5174504247638843, 0.29536587950758275, 12.762245750758076, 1.4412778801167454, 0.2805391871314324, 12.12161016992937, 1.368929023191677, 0.26645676084039477, 11.513133031700733, 1.3002119136003982, 0.2530812401773028, 10.935200055720887, 1.2349442459236248, 0.2403771400945878, 10.3862779948243, 1.1729528660576356, 0.22831075681300178, 9.864910567350384, 1.11407331183914, 0.21685007840601758, 9.369714593650976, 1.0581493767297228, 0.20596469987268715, 8.899376326536332, 1.0050326954023387, 0.19562574247364856, 8.452647965924314, 0.9545823501304124, 0.1858057771162812, 8.028344348446266, 0.9066644969353114, 0.17647875158575127, 7.62533980322708, 0.8611520105003578, 0.16761992142889215, 7.242565165497944, 0.8179241469093488, 0.1592057843075566, 6.879004940118887, 0.7768662233148302, 0.15121401764728032, 6.533694607486025, 0.7378693136862928, 0.14362341941584025, 6.205718064676107, 0.7008299598311127, 0.13641385187459415, 5.894205195039756, 0.6656498969215817, 0.129566188153374},
		'{-7.9971601676765065, -0.9647932237871281, 0.0674678376172424, -7.53640548355608, -1.0313925870870613, 0.049983942051968974, -7.042771240403503, -1.0868870463225866, 0.03301699880865099, -6.521623522189, -1.1314273786914566, 0.016667539808786005, -5.978260770751318, -1.1652385878824592, 0.0010263583421250763, -5.417877613529985, -1.188614440255397, -0.013825673700655287, -4.8455313103114905, -1.2019117652081905, -0.027817705098760373, -4.266110936455364, -1.2055445743624134, -0.04088892458692679, -3.684309393620352, -1.1999780527701942, -0.05298850408647032, -3.1045983132318247, -1.1857224735919805, -0.06407547018073582, -2.531205892977849, -1.1633270856458577, -0.07411850845148517, -1.9680976826378025, -1.1333740209153018, -0.08309570555959578, -1.4189603126635928, -1.0964722665542066, -0.09099423417017118, -0.8871881372648638, -1.0532517431767796, -0.09780998598971594, -0.37587274339591015, -1.0043575282963473, -0.103547158302657, 0.11220474191127638, -0.9504442607118933, -0.10821779946774397, 0.5745786309060368, -0.8921707584644062, -0.11184131886355088, 1.0091010421644866, -0.8301948797263012, -0.11444396675848531, 1.4139417707037965, -0.7651686526747791, -0.11605828952665566, 1.78758578934009, -0.6977336970615946, -0.11672256553911042}};
localparam real Fbi[0:2][0:59] = '{
	'{-2.7909677319823034, 1.1645589716088582, 0.19060596233437666, -3.3603178898584654, 1.0520184594053859, 0.19052933793233853, -3.8755368678013538, 0.9373449126732701, 0.18903196533224662, -4.3355298578492585, 0.8215044492173806, 0.18619741944199084, -4.7396707691325215, 0.7054226943956143, 0.18211501602510075, -5.087783031056338, 0.589979922753636, 0.1768788513948652, -5.380118013231764, 0.47600678626725107, 0.17058685528447062, -5.6173313449286635, 0.36428063124965954, 0.1633398633039268, -5.8004574181246475, 0.2555224014743813, 0.1552407149215018, -5.930882357334112, 0.1503941208060915, 0.14639338241404193, -6.010315736439308, 0.0494969446401462, 0.13690213572162893, -6.040761317838888, -0.046630234256533676, 0.12687074762212752, -6.024487082514156, -0.13751164332202986, 0.11640174311474336, -5.963994811231708, -0.22273497211670146, 0.10559569637302117, -5.861989467200935, -0.3019512222942703, 0.09455057810082401, -5.721348619237179, -0.37487409181022, 0.08336115560360488, -5.545092132000296, -0.44127892169979144, 0.07211844737531216, -5.336352336339004, -0.5010012355853093, 0.06090923350192322, -5.0983448783288265, -0.5539349035814157, 0.049815622698962225, -4.834340430399849, -0.6000299634619687, 0.03891467633524834},
	'{-8.958459938619613e-13, 2.0242635359008373e-14, 9.643826868290091e-15, -9.103308472692501e-13, 1.2512155407677278e-14, 7.852807227166043e-15, -9.211041253120783e-13, 5.506772714373422e-15, 6.217297157171153e-15, -9.285019541108567e-13, -8.268298269682301e-16, 4.7261972382432145e-15, -9.32836066726379e-13, -6.538443636357841e-15, 3.3691305267085744e-15, -9.343954051373796e-13, -1.1674554061510432e-14, 2.1363979903905273e-15, -9.334476228527553e-13, -1.6278546827448842e-14, 1.0189365973254915e-15, -9.302404940975976e-13, -2.0390902090185902e-14, 8.2799039720198e-18, -9.250032351662957e-13, -2.4049376818765866e-14, -9.034790024165938e-16, -9.179477432098616e-13, -2.728917618846588e-14, -1.7237223442930575e-15, -9.092697574171319e-13, -3.0143114628818584e-14, -2.459340406401403e-15, -8.991499472596516e-13, -3.264176713318623e-14, -3.116762322272564e-15, -8.877549321967428e-13, -3.481361140177142e-14, -3.701985009486355e-15, -8.75238236979681e-13, -3.668516135707408e-14, -4.220600361979052e-15, -8.617411864510661e-13, -3.828109253978835e-14, -4.677820801469937e-15, -8.473937435066098e-13, -3.9624359863872114e-14, -5.0785032842241965e-15, -8.323152936708476e-13, -4.073630818191976e-14, -5.427171853844682e-15, -8.166153795349887e-13, -4.163677608593021e-14, -5.7280388255720355e-15, -8.003943881135349e-13, -4.234419334400185e-14, -5.9850246826547555e-15, -7.837441939957622e-13, -4.287567235031996e-14, -6.201776760711041e-15},
	'{2.790967731983216, -1.164558971608878, -0.19060596233438637, 3.360317889859393, -1.0520184594053976, -0.19052933793234636, 3.8755368678022917, -0.9373449126732754, -0.18903196533225275, 4.335529857850204, -0.8215044492173792, -0.18619741944199542, 4.739670769133471, -0.7054226943956072, -0.18211501602510394, 5.087783031057288, -0.5899799227536234, -0.17687885139486717, 5.380118013232714, -0.4760067862672338, -0.17058685528447157, 5.617331344929609, -0.36428063124963816, -0.16333986330392686, 5.800457418125589, -0.25552240147435584, -0.1552407149215011, 5.930882357335045, -0.1503941208060623, -0.14639338241404057, 6.01031573644023, -0.04949694464011323, -0.13690213572162707, 6.040761317839798, 0.04663023425656987, -0.12687074762212525, 6.024487082515052, 0.13751164332206917, -0.1164017431147408, 5.963994811232588, 0.22273497211674398, -0.1055956963730184, 5.861989467201798, 0.3019512222943159, -0.09455057810082111, 5.721348619238023, 0.37487409181026843, -0.08336115560360194, 5.5450921320011215, 0.44127892169984273, -0.0721184473753092, 5.336352336339807, 0.5010012355853636, -0.06090923350192029, 5.098344878329605, 0.5539349035814728, -0.04981562269895935, 4.834340430400601, 0.6000299634620285, -0.03891467633524554}};
	localparam real hf[0:1199] = {0.030555386, 0.00018612405, -0.0001629881, 0.030435156, -5.2091487e-05, -0.0001618167, 0.030197391, -0.0002874397, -0.00015742924, 0.02984464, -0.0005178221, -0.00015012604, 0.029380444, -0.0007413086, -0.00014020878, 0.028809246, -0.000956142, -0.0001279783, 0.028136296, -0.0011607413, -0.00011373276, 0.027367568, -0.0013537037, -9.776573e-05, 0.026509656, -0.0015338041, -8.036446e-05, 0.025569687, -0.0016999954, -6.180824e-05, 0.024555236, -0.0018514054, -4.2366995e-05, 0.023474224, -0.0019873336, -2.229985e-05, 0.022334848, -0.002107248, -1.8539713e-06, 0.02114548, -0.0022107775, 1.8736506e-05, 0.019914603, -0.0022977078, 3.9251405e-05, 0.018650722, -0.002367973, 5.9485283e-05, 0.017362298, -0.002421649, 7.924808e-05, 0.01605768, -0.0024589433, 9.8365585e-05, 0.014745039, -0.002480188, 0.00011667984, 0.01343231, -0.0024858287, 0.00013404933, 0.012127141, -0.002476417, 0.00015034912, 0.01083684, -0.0024525977, 0.00016547077, 0.009568338, -0.0024151006, 0.00017932226, 0.008328148, -0.0023647302, 0.0001918277, 0.0071223313, -0.0023023542, 0.00020292701, 0.0059564738, -0.0022288947, 0.00021257541, 0.004835661, -0.0021453172, 0.00022074298, 0.003764464, -0.0020526215, 0.00022741394, 0.0027469255, -0.0019518309, 0.00023258604, 0.0017865527, -0.0018439849, 0.00023626979, 0.00088631624, -0.0017301285, 0.00023848764, 4.865055e-05, -0.0016113045, 0.00023927318, -0.00072454, -0.0014885457, 0.00023867021, -0.0014318712, -0.001362867, 0.00023673187, -0.002072466, -0.0012352585, 0.00023351966, -0.002645938, -0.0011066798, 0.00022910253, -0.003152372, -0.0009780528, 0.00022355597, -0.003592302, -0.00085025775, 0.00021696097, -0.0039666863, -0.0007241278, 0.00020940315, -0.004276882, -0.00060044543, 0.00020097184, -0.004524615, -0.00047993858, 0.00019175917, -0.004711952, -0.0003632781, 0.00018185917, -0.0048412695, -0.00025107525, 0.00017136698, -0.00491522, -0.00014388016, 0.00016037798, -0.004936704, -4.2180553e-05, 0.00014898712, -0.0049088323, 5.359881e-05, 0.00013728812, -0.0048348974, 0.00014309632, 0.00012537283, -0.0047183405, 0.00022601304, 0.00011333059, -0.004562718, 0.00030211205, 0.000101247715, -0.004371671, 0.00037121694, 8.9206915e-05, -0.0041488977, 0.00043321043, 7.7286866e-05, -0.003898119, 0.00048803218, 6.556179e-05, -0.003623056, 0.0005356765, 5.4101118e-05, -0.0033273993, 0.00057618966, 4.296917e-05, -0.0030147862, 0.0006096671, 3.2224943e-05, -0.002688776, 0.00063625025, 2.1921902e-05, -0.0023528298, 0.00065612316, 1.210784e-05, -0.0020102886, 0.0006695092, 2.8248041e-06, -0.0016643568, 0.00067666714, -5.890949e-06, -0.0013180855, 0.000677888, -1.4008946e-05, -0.00097435794, 0.00067349075, -2.1504444e-05, -0.000635878, 0.00066381897, -2.835834e-05, -0.00030515905, 0.0006492369, -3.4557037e-05, 1.5484078e-05, 0.00063012575, -4.009228e-05, 0.00032394167, 0.0006068802, -4.4960965e-05, 0.000618314, 0.0005799045, -4.9164897e-05, 0.00089691416, 0.00054960925, -5.2710555e-05, 0.0011582692, 0.0005164081, -5.560879e-05, 0.0014011202, 0.0004807144, -5.7874575e-05, 0.0016244196, 0.0004429382, -5.952664e-05, 0.0018273282, 0.00040348346, -6.058719e-05, 0.0020092104, 0.0003627453, -6.1081555e-05, 0.0021696282, 0.00032110757, -6.1037856e-05, 0.0023083335, 0.00027894066, -6.0486636e-05, 0.0024252608, 0.0002365993, -5.9460563e-05, 0.0025205174, 0.00019442089, -5.799403e-05, 0.0025943737, 0.00015272379, -5.6122874e-05, 0.0026472516, 0.00011180601, -5.3883978e-05, 0.0026797154, 7.194397e-05, -5.1315004e-05, 0.002692458, 3.3391636e-05, -4.8454043e-05, 0.00268629, -3.6202573e-06, -4.5339333e-05, 0.0026621271, -3.8884707e-05, -4.2008953e-05, 0.0026209771, -7.221876e-05, -3.8500562e-05, 0.0025639287, -0.00010346364, -3.4851157e-05, 0.002492138, -0.00013248467, -3.1096803e-05, 0.0024068162, -0.00015917102, -2.7272437e-05, 0.002309218, -0.00018343535, -2.3411669e-05, 0.0022006296, -0.00020521322, -1.954659e-05, 0.0020823576, -0.00022446235, -1.5707621e-05, 0.0019557173, -0.00024116186, -1.1923378e-05, 0.0018220227, -0.0002553113, -8.220541e-06, 0.0016825771, -0.0002669295, -4.623764e-06, 0.0015386626, -0.00027605367, -1.1556008e-06, 0.0013915325, -0.0002827379, 2.1635633e-06, 0.0012424025, -0.000287052, 5.315544e-06, 0.001092444, -0.00028908026, 8.284383e-06, 0.0009427772, -0.00028891992, 1.1056347e-05, 0.000794465, -0.00028667986, 1.3619921e-05, 0.0006485084, -0.00028247913, 1.5965776e-05, 0.00050584145, -0.00027644556, 1.8086721e-05, 0.00036732812, -0.0002687144, 1.9977653e-05, 0.00023375895, -0.00025942674, 2.1635487e-05, 0.000105848994, -0.00024872844, 2.3059069e-05, -1.5763893e-05, -0.0002367685, 2.4249082e-05, -0.0001305199, -0.00022369798, 2.5207959e-05, -0.00023793754, -0.00020966864, 2.5939764e-05, -0.0003376134, -0.00019483182, 2.6450076e-05, -0.00042922117, -0.00017933731, 2.6745873e-05, -0.00051251025, -0.00016333231, 2.6835407e-05, -0.0005873039, -0.00014696043, 2.6728076e-05, -0.0006534967, -0.00013036082, 2.643429e-05, -0.0007110519, -0.00011366732, 2.596535e-05, -0.0007599983, -9.70078e-05, 2.5333306e-05, -0.0008004264, -8.05034e-05, 2.455083e-05, -0.00083248515, -6.426804e-05, 2.36311e-05, -0.0008563774, -4.840788e-05, 2.258766e-05, -0.00087235606, -3.3020973e-05, 2.1434305e-05, -0.00088071957, -1.8196892e-05, 2.0184969e-05, -0.00088180724, -4.0165096e-06, 1.8853601e-05, -0.00087599485, 9.4481675e-06, 1.7454076e-05, -0.00086369005, 2.2134092e-05, 1.600008e-05, -0.0008453275, 3.398719e-05, 1.4505019e-05, -0.0008213646, 4.4962322e-05, 1.298194e-05, -0.0007922764, 5.502315e-05, 1.1443444e-05, -0.000758552, 6.4141976e-05, 9.901617e-06, -0.00072068936, 7.229951e-05, 8.367962e-06, -0.00067919167, 7.948459e-05, 6.8533486e-06, -0.0006345633, 8.569385e-05, 5.367956e-06, -0.0005873056, 9.093134e-05, 3.921237e-06, -0.000537914, 9.5208154e-05, 2.5218808e-06, -0.0004868739, 9.854194e-05, 1.1777888e-06, -0.0004346582, 0.00010095648, -1.0394647e-07, -0.00038172395, 0.000102481186, -1.3170527e-06, -0.00032851, 0.00010315059, -2.4560836e-06, -0.0002754347, 0.00010300382, -3.516418e-06, -0.0002228936, 0.000102084094, -4.4942517e-06, -0.00017125793, 0.000100438185, -5.3865865e-06, -0.000120872864, 9.811589e-05, -6.19121e-06, -7.205645e-05, 9.5169475e-05, -6.9066728e-06, -2.5098529e-05, 9.165322e-05, -7.5322623e-06, 1.9739968e-05, 8.762287e-05, -8.067968e-06, 6.222746e-05, 8.313514e-05, -8.514448e-06, 0.00010216197, 7.824727e-05, -8.872992e-06, 0.0001393711, 7.301654e-05, -9.145473e-06, 0.00017371179, 6.749988e-05, -9.3343115e-06, 0.00020506994, 6.1753424e-05, -9.442427e-06, 0.0002333597, 5.583216e-05, -9.473187e-06, 0.0002585227, 4.9789553e-05, -9.430366e-06, 0.00028052714, 4.3677246e-05, -9.3180915e-06, 0.0002993665, 3.754476e-05, -9.140798e-06, 0.00031505854, 3.1439224e-05, -8.903177e-06, 0.00032764368, 2.5405157e-05, -8.610128e-06, 0.00033718365, 1.9484261e-05, -8.266716e-06, 0.00034375995, 1.371526e-05, -7.878119e-06, 0.00034747223, 8.133754e-06, -7.4495883e-06, 0.00034843653, 2.772119e-06, -6.9864045e-06, 0.00034678367, -2.3405717e-06, -6.493835e-06, 0.00034265747, -7.1785967e-06, -5.977097e-06, 0.00033621298, -1.1719608e-05, -5.4413213e-06, 0.00032761483, -1.5944624e-05, -4.8915176e-06, 0.00031703542, -1.9838002e-05, -4.332543e-06, 0.00030465322, -2.3387383e-05, -3.7690756e-06, 0.00029065125, -2.6583617e-05, -3.2055857e-06, 0.00027521534, -2.9420667e-05, -2.6463154e-06, 0.00025853264, -3.18955e-05, -2.0952575e-06, 0.0002407902, -3.4007942e-05, -1.5561386e-06, 0.00022217346, -3.5760553e-05, -1.0324053e-06, 0.00020286506, -3.7158454e-05, -5.272122e-07, 0.00018304354, -3.8209168e-05, -4.3413344e-08, 0.00016288225, -3.8922426e-05, 4.1644353e-07, 0.00014254828, -3.9309998e-05, 8.5012056e-07, 0.00012220157, -3.9385497e-05, 1.2556906e-06, 0.00010199404, -3.9164173e-05, 1.6315356e-06, 8.206888e-05, -3.8662725e-05, 1.9763434e-06, 6.2559906e-05, -3.7899106e-05, 2.2891013e-06, 4.3591048e-05, -3.6892307e-05, 2.5690888e-06, 2.5275926e-05, -3.566218e-05, 2.8158674e-06, 7.717512e-06, -3.4229237e-05, 3.0292708e-06, -8.992086e-06, -3.2614473e-05, 3.209391e-06, -2.477177e-05, -3.083916e-05, 3.3565643e-06, -3.95515e-05, -2.8924704e-05, 3.4713576e-06, -5.327225e-05, -2.6892454e-05, 3.554551e-06, -6.5885884e-05, -2.4763562e-05, 3.6071226e-06, -7.735499e-05, -2.2558823e-05, 3.630229e-06, -8.7652574e-05, -2.0298543e-05, 3.6251893e-06, -9.676176e-05, -1.800241e-05, 3.593466e-06, -0.000104675404, -1.5689382e-05, 3.536648e-06, -0.00011139564, -1.3377577e-05, 3.45643e-06, -0.00011693339, -1.1084184e-05, 3.3545969e-06, -0.00012130786, -8.825379e-06, 3.2330036e-06, -0.00012454593, -6.616259e-06, 3.0935591e-06, -0.0001266816, -4.4707804e-06, 2.9382095e-06, -0.0001277554, -2.4017152e-06, 2.7689205e-06, -0.00012781366, -4.206141e-07, 2.5876618e-06, -0.00012690797, 1.4622167e-06, 2.3963933e-06, -0.00012509448, 3.2377293e-06, 2.1970495e-06, -0.00012243325, 4.8981383e-06, 1.9915278e-06, -0.00011898759, 6.4369146e-06, 1.7816747e-06, -0.000114823466, 7.848769e-06, 1.5692755e-06, -0.00011000883, 9.129632e-06, 1.3560439e-06, -0.00010461302, 1.0276617e-05, 1.1436125e-06, -9.870619e-05, 1.1287986e-05, 9.3352514e-07, -9.235872e-05, 1.2163104e-05, 7.2722963e-07, -8.5640706e-05, 1.2902383e-05, 5.260719e-07, -7.862142e-05, 1.3507232e-05, 3.3129098e-07, -7.136885e-05, 1.3979992e-05, 1.4401532e-07, -6.394926e-05, 1.432387e-05, -3.474011e-08, -5.6426783e-05, 1.4542874e-05, -2.0407558e-07, -4.8863043e-05, 1.4641741e-05, -3.6320748e-07, -4.131683e-05, 1.4625863e-05, -5.1146833e-07, -3.3843797e-05, 1.4501216e-05, -6.4830573e-07, -2.649621e-05, 1.4274286e-05, -7.732808e-07, -1.932273e-05, 1.3951988e-05, -8.8606555e-07, -1.236823e-05, 1.3541601e-05, -9.864398e-07, -5.6736553e-06, 1.30506905e-05, -1.0742872e-06, 7.240838e-07, 1.24870385e-05, -1.149591e-06, 6.7921815e-06, 1.1858574e-05, -1.2124287e-06, 1.2501972e-05, 1.1173305e-05, -1.2629675e-06, 1.7828936e-05, 1.04392575e-05, -1.3014576e-06, 2.2752663e-05, 9.664412e-06, -1.3282264e-06, 2.7256812e-05, 8.856648e-06, -1.3436725e-06, 3.1329004e-05, 8.023688e-06, -1.3482585e-06, 3.4960736e-05, 7.1730506e-06, -1.3425046e-06, 3.814722e-05, 6.312003e-06, -1.326982e-06, 4.0887262e-05, 5.447519e-06, -1.3023055e-06, 4.3183056e-05, 4.5862425e-06, -1.2691271e-06, 4.504001e-05, 3.7344562e-06, -1.228129e-06, 4.646655e-05, 2.8980496e-06, -1.1800173e-06, 4.7473888e-05, 2.0824982e-06, -1.125515e-06, 4.80758e-05, 1.2928417e-06, -1.0653561e-06, 4.8288395e-05, 5.336698e-07, -1.0002794e-06, 4.8129874e-05, -1.9089032e-07, -9.310231e-07, 4.762029e-05, -8.7718036e-07, -8.583185e-07, 4.6781304e-05, -1.5220149e-06, -7.828858e-07, 4.563593e-05, -2.1226808e-06, -7.054287e-07, 4.420831e-05, -2.676934e-06, -6.266301e-07, 4.2523465e-05, -3.1829911e-06, -5.4714826e-07, 4.060707e-05, -3.6395209e-06, -4.6761284e-07, 3.8485214e-05, -4.0456302e-06, -3.886219e-07, 3.6184207e-05, -4.400849e-06, -3.1073893e-07, 3.3730354e-05, -4.70511e-06, -2.3449027e-07, 3.1149768e-05, -4.958733e-06, -1.6036336e-07, 2.8468174e-05, -5.162399e-06, -8.880481e-08, 2.5710748e-05, -5.317127e-06, -2.0219318e-08, 2.290195e-05, -5.4242523e-06, 4.5031335e-08, 2.0065378e-05, -5.4853967e-06, 1.0662873e-07, 1.7223641e-05, -5.502444e-06, 1.6429802e-07, 1.439823e-05, -5.477511e-06, 2.1780772e-07, 1.16094225e-05, -5.4129214e-06, 2.6696932e-07, 8.876192e-06, -5.3111767e-06, 3.116364e-07, 6.216127e-06, -5.1749294e-06, 3.517036e-07, 3.6453769e-06, -5.0069543e-06, 3.8710536e-07, 1.178599e-06, -4.810123e-06, 4.178144e-07, -1.1710715e-06, -4.5873753e-06, 4.438399e-07, -3.392044e-06, -4.3416962e-06, 4.6522558e-07, -5.47428e-06, -4.07609e-06, 4.8204765e-07, -7.4092886e-06, -3.7935565e-06, 4.9441263e-07, -9.190113e-06, -3.4970699e-06, 5.024549e-07, -1.0811303e-05, -3.1895568e-06, 5.063343e-07, -1.2268877e-05, -2.8738775e-06, 5.0623373e-07, -1.3560282e-05, -2.5528077e-06, 5.0235656e-07, -1.4684335e-05, -2.2290217e-06, 4.949239e-07, -1.5641166e-05, -1.9050784e-06, 4.8417235e-07, -1.6432148e-05, -1.5834072e-06, 4.7035118e-07, -1.7059821e-05, -1.2662967e-06, 4.5372e-07, -1.752782e-05, -9.558853e-07, 4.345462e-07, -1.7840786e-05, -6.541521e-07, 4.1310247e-07, -1.8004284e-05, -3.6291038e-07, 3.8966473e-07, -1.8024713e-05, -8.380295e-08, 3.6450967e-07, -1.7909213e-05, 1.8170195e-07, 3.3791275e-07, -1.7665578e-05, 4.3231256e-07, 3.101462e-07, -1.7302164e-05, 6.669142e-07, 2.814771e-07, -1.6827795e-05, 8.8456875e-07, 2.521657e-07, -1.6251674e-05, 1.0845125e-06, 2.2246381e-07, -1.5583299e-05, 1.2661532e-06, 1.9261331e-07, -1.4832369e-05, 1.4290653e-06, 1.6284491e-07, -1.4008711e-05, 1.5729852e-06, 1.3337691e-07, -1.3122193e-05, 1.6978047e-06, 1.044143e-07, -1.2182649e-05, 1.8035638e-06, 7.614779e-08, -1.1199809e-05, 1.8904433e-06, 4.8753233e-08, -1.018323e-05, 1.9587553e-06, 2.2390962e-08, -9.142238e-06, 2.0089356e-06, -2.7945448e-09, -8.085861e-06, 2.0415325e-06, -2.6674979e-08, -7.0227857e-06, 2.0571986e-06, -4.913832e-08, -5.961305e-06, 2.0566797e-06, -7.0088845e-08, -4.909277e-06, 2.040804e-06, -8.944703e-08, -3.8740886e-06, 2.010473e-06, -1.07149276e-07, -2.862625e-06, 1.9666502e-06, -1.2314764e-07, -1.8812433e-06, 1.9103509e-06, -1.3740934e-07, -9.357506e-07, 1.8426315e-06, -1.4991626e-07, -3.139061e-08, 1.7645806e-06, -1.606643e-07, 8.271681e-07, 1.6773082e-06, -1.6966274e-07, 1.6358373e-06, 1.5819369e-06, -1.7693347e-07, 2.3911102e-06, 1.4795925e-06, -1.8251016e-07, 3.090058e-06, 1.3713956e-06, -1.8643746e-07, 3.7303223e-06, 1.2584537e-06, -1.8877006e-07, 4.3101036e-06, 1.141853e-06, -1.8957176e-07, 4.8281468e-06, 1.022652e-06, -1.8891463e-07, 5.2837217e-06, 9.018745e-07, -1.868779e-07, 5.676604e-06, 7.8050414e-07, -1.835471e-07, 6.0070474e-06, 6.5947864e-07, -1.790131e-07, 6.2757613e-06, 5.396855e-07, -1.7337112e-07, 6.48388e-06, 4.2195788e-07, -1.667198e-07, 6.632934e-06, 3.0707082e-07, -1.5916032e-07, 6.7248156e-06, 1.9573879e-07, -1.507955e-07, 6.7617502e-06, 8.8613255e-08, -1.4172892e-07, 6.74626e-06, -1.3719013e-08, -1.3206414e-07, 6.6811303e-06, -1.1073694e-07, -1.2190394e-07, 6.5693766e-06, -2.0198576e-07, -1.1134951e-07, 6.4142087e-06, -2.87077e-07, -1.0049989e-07, 6.218998e-06, -3.65688e-07, -8.9451255e-08, 5.987243e-06, -4.375611e-07, -7.8296374e-08, 5.7225384e-06, -5.02502e-07, -6.712408e-08, 5.428541e-06, -5.603783e-07, -5.6018806e-08, 5.1089405e-06, -6.1111695e-07, -4.506019e-08, 4.767431e-06, -6.5470226e-07, -3.4322714e-08, 4.407682e-06, -6.9117266e-07, -2.3875408e-08, 4.033311e-06, -7.2061783e-07, -1.3781621e-08, 3.647863e-06, -7.4317546e-07, -4.0988235e-09, 3.254783e-06, -7.590277e-07, 5.1215094e-09, 2.857399e-06, -7.683977e-07, 1.3833986e-08, 2.4589015e-06, -7.7154544e-07, 2.1999325e-08, 2.0623258e-06, -7.687644e-07, 2.9584337e-08, 1.6705397e-06, -7.6037736e-07, 3.656186e-08, 1.2862281e-06, -7.4673255e-07, 4.291067e-08, 9.118834e-07, -7.2819995e-07, 4.861531e-08, 5.497967e-07, -7.05167e-07, 5.3665936e-08, 2.0205074e-07, -6.780352e-07, 5.8058095e-08, -1.2948513e-07, -6.4721615e-07, 6.1792484e-08, -4.4315803e-07, -6.131282e-07, 6.487469e-08, -7.3753273e-07, -5.761927e-07, 6.731488e-08, -1.0113915e-06, -5.3683084e-07, 6.9127516e-08, -1.263732e-06, -4.954606e-07, 7.0331e-08, -1.4937638e-06, -4.524936e-07, 7.0947365e-08, -1.7009036e-06, -4.083324e-07, 7.1001914e-08, -1.884769e-06, -3.6336806e-07, 7.052285e-08, -2.045171e-06, -3.1797768e-07, 6.9540945e-08, -2.1821056e-06, -2.7252236e-07, 6.808914e-08, -2.2957447e-06, -2.2734525e-07, 6.620224e-08, -2.3864256e-06, -1.8277e-07, 6.39165e-08, -2.4546398e-06, -1.3909921e-07, 6.126935e-08, -2.501022e-06, -9.6613356e-08, 5.8298966e-08, -2.526338e-06, -5.556973e-08, 5.504404e-08, -2.5314714e-06, -1.620174e-08, 5.1543402e-08, -2.5174122e-06, 2.1281616e-08, 4.7835737e-08, -2.4852436e-06, 5.6696084e-08, 4.3959314e-08, -2.4361286e-06, 8.988227e-08, 3.9951715e-08, -2.371298e-06, 1.2070555e-07, 3.5849588e-08, -2.2920374e-06, 1.4905585e-07, 3.168842e-08, -2.1996743e-06, 1.7484716e-07, 2.7502324e-08, -2.0955672e-06, 1.98017e-07, 2.3323878e-08, -1.981093e-06, 2.185257e-07, 1.918393e-08, -1.8576355e-06, 2.3635546e-07, 1.5111471e-08, -1.7265759e-06, 2.5150945e-07, 1.1133516e-08, -1.5892814e-06, 2.640107e-07, 7.274993e-09, -1.4470963e-06, 2.7390087e-07, 3.5586671e-09, -1.301333e-06, 2.81239e-07, 5.0811855e-12, -1.1532638e-06, 2.8610032e-07, -3.3674854e-09, -1.0041133e-06, 2.8857457e-07, -6.5430377e-09, -8.55052e-07, 2.887649e-07, -9.507868e-09, -7.0718994e-07, 2.8678627e-07, -1.22505455e-08, -5.6157165e-07, 2.8276395e-07, -1.4761879e-08, -4.1917178e-07, 2.7683214e-07, -1.7034878e-08, -2.808912e-07, 2.6913244e-07, -1.9064688e-08, -1.4755398e-07, 2.5981257e-07, -2.0848521e-08, -1.9905396e-08, 2.4902468e-07, -2.2385573e-08, 1.01389844e-07, 2.3692427e-07, -2.367692e-08, 2.1574841e-07, 2.2366866e-07, -2.4725427e-08, 3.2266857e-07, 2.0941584e-07, -2.5535627e-08, 4.217297e-07, 1.9432319e-07, -2.6113598e-08, 5.125915e-07, 1.7854634e-07, -2.6466855e-08, 5.949922e-07, 1.6223812e-07, -2.6604202e-08, 6.687466e-07, 1.4554755e-07, -2.6535611e-08, 7.3374383e-07, 1.286189e-07, -2.627209e-08, 7.8994384e-07, 1.1159089e-07, -2.5825539e-08, 8.373746e-07, 9.459591e-08, -2.5208621e-08, 8.761282e-07, 7.775936e-08, -2.4434629e-08, 9.0635683e-07, 6.119905e-08, -2.3517352e-08, 9.282688e-07, 4.502475e-08, -2.247095e-08, 9.421238e-07, 2.933773e-08, -2.1309825e-08, 9.4822883e-07, 1.4230468e-08, -2.0048505e-08, 9.4693297e-07, -2.1360864e-10, -1.8701526e-08, 9.386229e-07, -1.392028e-08, -1.7283321e-08, 9.237181e-07, -2.6824623e-08, -1.5808128e-08, 9.02666e-07, -3.8871015e-08, -1.4289878e-08, 8.759371e-07, -5.0013092e-08, -1.2742118e-08, 8.440204e-07, -6.021361e-08, -1.11779235e-08, 8.07419e-07, -6.9444255e-08, -9.60983e-09, 7.6664503e-07, -7.768542e-08, -8.049761e-09, 7.2221604e-07, -8.4925894e-08, -6.508972e-09, 6.7465044e-07, -9.1162505e-08, -4.9980033e-09, 6.244636e-07, -9.6399766e-08, -3.5266332e-09, 5.7216437e-07, -1.0064943e-07, -2.1038469e-09, 5.182514e-07, -1.0393002e-07, -7.378082e-10, 4.6320997e-07, -1.06266384e-07, 5.6415944e-10, 4.075092e-07, -1.0768915e-07, 1.7955847e-09, 3.515991e-07, -1.0823422e-07, 2.9508531e-09, 2.9590845e-07, -1.07942235e-07, 4.0252064e-09, 2.408424e-07, -1.0685802e-07, 5.0147326e-09, 1.8678092e-07, -1.0503003e-07, 5.9163545e-09};
	localparam real hb[0:1199] = {0.030555386, 0.00042473868, -0.00016067282, 0.030435156, 0.00066057424, -0.00015489412, 0.030197391, 0.0008911913, -0.00014596741, 0.02984464, 0.0011145421, -0.00013423445, 0.029380444, 0.0013287675, -0.000120034856, 0.028809246, 0.0015321989, -0.000103703904, 0.028136296, 0.0017233604, -8.557052e-05, 0.027367568, 0.0019009683, -6.595545e-05, 0.026509656, 0.0020639296, -4.516946e-05, 0.025569687, 0.0022113395, -2.3511817e-05, 0.024555236, 0.0023424772, -1.2688207e-06, 0.023474224, 0.0024568012, 2.1287447e-05, 0.022334848, 0.0025539424, 4.3900236e-05, 0.02114548, 0.0026336978, 6.632907e-05, 0.019914603, 0.0026960226, 8.835055e-05, 0.018650722, 0.002741021, 0.00010975895, 0.017362298, 0.002768938, 0.00013036674, 0.01605768, 0.0027801483, 0.00015000484, 0.014745039, 0.002775147, 0.00016852286, 0.01343231, 0.0027545395, 0.0001857891, 0.012127141, 0.002719029, 0.00020169046, 0.01083684, 0.0026694075, 0.00021613219, 0.009568338, 0.0026065432, 0.00022903756, 0.008328148, 0.0025313706, 0.0002403474, 0.0071223313, 0.002444879, 0.00025001957, 0.0059564738, 0.0023481022, 0.00025802825, 0.004835661, 0.0022421074, 0.0002643632, 0.003764464, 0.0021279857, 0.000269029, 0.0027469255, 0.002006842, 0.00027204418, 0.0017865527, 0.0018797856, 0.00027344024, 0.00088631624, 0.0017479206, 0.00027326067, 4.865055e-05, 0.0016123392, 0.00027155995, -0.00072454, 0.0014741119, 0.00026840257, -0.0014318712, 0.0013342815, 0.00026386188, -0.002072466, 0.001193856, 0.00025801905, -0.002645938, 0.0010538022, 0.00025096207, -0.003152372, 0.0009150408, 0.00024278458, -0.003592302, 0.00077844126, 0.00023358493, -0.0039666863, 0.0006448177, 0.00022346506, -0.004276882, 0.0005149255, 0.00021252957, -0.004524615, 0.00038945812, 0.00020088472, -0.004711952, 0.00026904506, 0.00018863752, -0.0048412695, 0.00015425023, 0.00017589486, -0.00491522, 4.5570643e-05, 0.00016276263, -0.004936704, -5.6563887e-05, 0.00014934501, -0.0049088323, -0.00015179084, 0.00013574367, -0.0048348974, -0.00023981437, 0.00012205715, -0.0047183405, -0.00032040442, 0.000108380234, -0.004562718, -0.00039339505, 9.480342e-05, -0.004371671, -0.00045868277, 8.141238e-05, -0.0041488977, -0.0005162242, 6.82876e-05, -0.003898119, -0.0005660334, 5.5503962e-05, -0.003623056, -0.00060817914, 4.3130498e-05, -0.0033273993, -0.00064278144, 3.123009e-05, -0.0030147862, -0.0006700085, 1.9859337e-05, -0.002688776, -0.00069007295, 9.068396e-06, -0.0023528298, -0.0007032281, -1.0990615e-06, -0.0020102886, -0.000709764, -1.060588e-05, -0.0016643568, -0.00071000383, -1.9421377e-05, -0.0013180855, -0.0007042993, -2.7521268e-05, -0.00097435794, -0.0006930272, -3.488753e-05, -0.000635878, -0.0006765853, -4.150824e-05, -0.00030515905, -0.000655388, -4.737736e-05, 1.5484078e-05, -0.0006298628, -5.2494524e-05, 0.00032394167, -0.0006004467, -5.6864723e-05, 0.000618314, -0.0005675819, -6.049804e-05, 0.00089691416, -0.00053171284, -6.340932e-05, 0.0011582692, -0.00049328257, -6.561782e-05, 0.0014011202, -0.00045272967, -6.7146866e-05, 0.0016244196, -0.00041048517, -6.8023466e-05, 0.0018273282, -0.0003669698, -6.827794e-05, 0.0020092104, -0.00032259143, -6.794353e-05, 0.0021696282, -0.0002777427, -6.705603e-05, 0.0023083335, -0.00023279902, -6.565337e-05, 0.0024252608, -0.0001881164, -6.377523e-05, 0.0025205174, -0.00014403016, -6.146269e-05, 0.0025943737, -0.00010085325, -5.8757854e-05, 0.0026472516, -5.887523e-05, -5.5703462e-05, 0.0026797154, -1.8361296e-05, -5.234257e-05, 0.002692458, 2.044845e-05, -4.871821e-05, 0.00268629, 5.7339465e-05, -4.487308e-05, 0.0026621271, 9.2123046e-05, -4.0849245e-05, 0.0026209771, 0.00012463638, -3.6687852e-05, 0.0025639287, 0.00015474246, -3.2428892e-05, 0.002492138, 0.0001823297, -2.8110948e-05, 0.0024068162, 0.00020731153, -2.3770992e-05, 0.002309218, 0.00022962567, -1.9444191e-05, 0.0022006296, 0.0002492334, -1.5163747e-05, 0.0020823576, 0.00026611856, -1.0960741e-05, 0.0019557173, 0.0002802866, -6.8640243e-06, 0.0018220227, 0.00029176328, -2.9001133e-06, 0.0016825771, 0.00030059362, 9.068854e-07, 0.0015386626, 0.00030684032, 4.535327e-06, 0.0013915325, 0.00031058263, 7.966065e-06, 0.0012424025, 0.00031191471, 1.118246e-05, 0.001092444, 0.00031094422, 1.41703795e-05, 0.0009427772, 0.00030779082, 1.6918166e-05, 0.000794465, 0.00030258464, 1.9416602e-05, 0.0006485084, 0.0002954648, 2.1658849e-05, 0.00050584145, 0.00028657776, 2.3640374e-05, 0.00036732812, 0.00027607608, 2.5358868e-05, 0.00023375895, 0.0002641167, 2.6814143e-05, 0.000105848994, 0.00025085977, 2.8008028e-05, -1.5763893e-05, 0.00023646705, 2.8944247e-05, -0.0001305199, 0.0002211008, 2.9628292e-05, -0.00023793754, 0.00020492243, 3.00673e-05, -0.0003376134, 0.00018809135, 3.0269897e-05, -0.00042922117, 0.00017076389, 3.0246076e-05, -0.00051251025, 0.00015309226, 3.000703e-05, -0.0005873039, 0.00013522363, 2.9565026e-05, -0.0006534967, 0.00011729925, 2.8933244e-05, -0.0007110519, 9.9453726e-05, 2.8125638e-05, -0.0007599983, 8.181434e-05, 2.7156782e-05, -0.0008004264, 6.450043e-05, 2.604174e-05, -0.00083248515, 4.7622954e-05, 2.479592e-05, -0.0008563774, 3.1284024e-05, 2.3434939e-05, -0.00087235606, 1.557663e-05, 2.1974502e-05, -0.00088071957, 5.8439167e-07, 2.0430272e-05, -0.00088180724, -1.3618604e-05, 1.8817758e-05, -0.00087599485, -2.6967859e-05, 1.7152202e-05, -0.00086369005, -3.9408475e-05, 1.5448486e-05, -0.0008453275, -5.089507e-05, 1.372103e-05, -0.0008213646, -6.1391635e-05, 1.1983708e-05, -0.0007922764, -7.087135e-05, 1.0249777e-05, -0.000758552, -7.931628e-05, 8.531804e-06, -0.00072068936, -8.671711e-05, 6.841608e-06, -0.00067919167, -9.307273e-05, 5.190208e-06, -0.0006345633, -9.838985e-05, 3.5877833e-06, -0.0005873056, -0.00010268257, 2.043637e-06, -0.000537914, -0.00010597187, 5.661719e-07, -0.0004868739, -0.00010828512, -8.37127e-07, -0.0004346582, -0.000109655564, -2.1597023e-06, -0.00038172395, -0.00011012174, -3.3959263e-06, -0.00032851, -0.00010972696, -4.541096e-06, -0.0002754347, -0.00010851874, -5.5914225e-06, -0.0002228936, -0.00010654821, -6.5440113e-06, -0.00017125793, -0.00010386954, -7.396841e-06, -0.000120872864, -0.00010053946, -8.148731e-06, -7.205645e-05, -9.66166e-05, -8.799312e-06, -2.5098529e-05, -9.2161026e-05, -9.348984e-06, 1.9739968e-05, -8.7233704e-05, -9.798878e-06, 6.222746e-05, -8.1895996e-05, -1.0150804e-05, 0.00010216197, -7.620917e-05, -1.0407213e-05, 0.0001393711, -7.023398e-05, -1.0571139e-05, 0.00017371179, -6.403021e-05, -1.0646147e-05, 0.00020506994, -5.765627e-05, -1.0636282e-05, 0.0002333597, -5.116887e-05, -1.0546015e-05, 0.0002585227, -4.462266e-05, -1.0380185e-05, 0.00028052714, -3.806991e-05, -1.0143948e-05, 0.0002993665, -3.1560274e-05, -9.84272e-06, 0.00031505854, -2.5140533e-05, -9.482121e-06, 0.00032764368, -1.88544e-05, -9.0679305e-06, 0.00033718365, -1.2742346e-05, -8.606027e-06, 0.00034375995, -6.841464e-06, -8.102347e-06, 0.00034747223, -1.1853657e-06, -7.5628327e-06, 0.00034843653, 4.195892e-06, -6.9933894e-06, 0.00034678367, 9.27585e-06, -6.399843e-06, 0.00034265747, 1.4031661e-05, -5.7879006e-06, 0.00033621298, 1.8444078e-05, -5.1631146e-06, 0.00032761483, 2.2497408e-05, -4.5308484e-06, 0.00031703542, 2.6179458e-05, -3.8962453e-06, 0.00030465322, 2.9481436e-05, -3.264203e-06, 0.00029065125, 3.2397853e-05, -2.6393498e-06, 0.00027521534, 3.4926386e-05, -2.0260213e-06, 0.00025853264, 3.706774e-05, -1.4282452e-06, 0.0002407902, 3.8825492e-05, -8.4972646e-07, 0.00022217346, 4.020591e-05, -2.9383557e-07, 0.00020286506, 4.1217758e-05, 2.3639892e-07, 0.00018304354, 4.1872132e-05, 7.3829597e-07, 0.00016288225, 4.218224e-05, 1.2095242e-06, 0.00014254828, 4.216319e-05, 1.6481011e-06, 0.00012220157, 4.1831787e-05, 2.052391e-06, 0.00010199404, 4.1206327e-05, 2.4210985e-06, 8.206888e-05, 4.0306375e-05, 2.753261e-06, 6.2559906e-05, 3.9152554e-05, 3.0482397e-06, 4.3591048e-05, 3.7766342e-05, 3.305707e-06, 2.5275926e-05, 3.6169862e-05, 3.5256328e-06, 7.717512e-06, 3.4385692e-05, 3.7082707e-06, -8.992086e-06, 3.2436656e-05, 3.8541407e-06, -2.477177e-05, 3.0345662e-05, 3.964012e-06, -3.95515e-05, 2.8135513e-05, 4.038884e-06, -5.327225e-05, 2.5828742e-05, 4.079968e-06, -6.5885884e-05, 2.3447463e-05, 4.0886675e-06, -7.735499e-05, 2.101322e-05, 4.0665554e-06, -8.7652574e-05, 1.8546863e-05, 4.0153573e-06, -9.676176e-05, 1.6068418e-05, 3.936927e-06, -0.000104675404, 1.3596983e-05, 3.83323e-06, -0.00011139564, 1.115064e-05, 3.7063194e-06, -0.00011693339, 8.746357e-06, 3.558319e-06, -0.00012130786, 6.399928e-06, 3.3914012e-06, -0.00012454593, 4.1259145e-06, 3.207771e-06, -0.0001266816, 1.937592e-06, 3.0096453e-06, -0.0001277554, -1.5307594e-07, 2.7992373e-06, -0.00012781366, -2.1354654e-06, 2.5787397e-06, -0.00012690797, -4.0003006e-06, 2.350309e-06, -0.00012509448, -5.739656e-06, 2.1160513e-06, -0.00012243325, -7.3469473e-06, 1.87801e-06, -0.00011898759, -8.816911e-06, 1.6381523e-06, -0.000114823466, -1.0145576e-05, 1.3983592e-06, -0.00011000883, -1.1330232e-05, 1.1604159e-06, -0.00010461302, -1.236938e-05, 9.2600254e-07, -9.870619e-05, -1.3262684e-05, 6.96688e-07, -9.235872e-05, -1.4010915e-05, 4.739231e-07, -8.5640706e-05, -1.4615889e-05, 2.59036e-07, -7.862142e-05, -1.50804e-05, 5.322848e-08, -7.136885e-05, -1.5408146e-05, -1.4242659e-07, -6.394926e-05, -1.5603664e-05, -3.2698674e-07, -5.6426783e-05, -1.5672242e-05, -4.996403e-07, -4.8863043e-05, -1.5619851e-05, -6.5970585e-07, -4.131683e-05, -1.5453059e-05, -8.066306e-07, -3.3843797e-05, -1.5178954e-05, -9.399882e-07, -2.649621e-05, -1.4805067e-05, -1.059475e-06, -1.932273e-05, -1.4339289e-05, -1.1649067e-06, -1.236823e-05, -1.3789796e-05, -1.2562134e-06, -5.6736553e-06, -1.3164972e-05, -1.333434e-06, 7.240838e-07, -1.247334e-05, -1.3967109e-06, 6.7921815e-06, -1.1723481e-05, -1.4462831e-06, 1.2501972e-05, -1.0923982e-05, -1.4824802e-06, 1.7828936e-05, -1.0083357e-05, -1.5057145e-06, 2.2752663e-05, -9.209995e-06, -1.5164744e-06, 2.7256812e-05, -8.312103e-06, -1.5153166e-06, 3.1329004e-05, -7.3976535e-06, -1.5028584e-06, 3.4960736e-05, -6.4743335e-06, -1.47977e-06, 3.814722e-05, -5.5495066e-06, -1.4467672e-06, 4.0887262e-05, -4.6301716e-06, -1.4046028e-06, 4.3183056e-05, -3.722929e-06, -1.3540604e-06, 4.504001e-05, -2.8339527e-06, -1.2959457e-06, 4.646655e-05, -1.968965e-06, -1.2310801e-06, 4.7473888e-05, -1.1332174e-06, -1.1602938e-06, 4.80758e-05, -3.314743e-07, -1.0844185e-06, 4.8288395e-05, 4.3199668e-07, -1.004282e-06, 4.8129874e-05, 1.1534319e-06, -9.2070127e-07, 4.762029e-05, 1.8295738e-06, -8.344777e-07, 4.6781304e-05, 2.45767e-06, -7.4639155e-07, 4.563593e-05, 3.0354677e-06, -6.57197e-07, 4.420831e-05, 3.5612047e-06, -5.6761826e-07, 4.2523465e-05, 4.033599e-06, -4.783454e-07, 4.060707e-05, 4.451832e-06, -3.9003106e-07, 3.8485214e-05, 4.8155325e-06, -3.0328738e-07, 3.6184207e-05, 5.124756e-06, -2.1868355e-07, 3.3730354e-05, 5.379963e-06, -1.3674376e-07, 3.1149768e-05, 5.5819937e-06, -5.794553e-08, 2.8468174e-05, 5.732044e-06, 1.7281472e-08, 2.5710748e-05, 5.8316373e-06, 8.855619e-08, 2.290195e-05, 5.882597e-06, 1.5554656e-07, 2.0065378e-05, 5.8870182e-06, 2.1796949e-07, 1.7223641e-05, 5.8472356e-06, 2.7559048e-07, 1.439823e-05, 5.7657967e-06, 3.282229e-07, 1.16094225e-05, 5.6454305e-06, 3.7572698e-07, 8.876192e-06, 5.489019e-06, 4.1800843e-07, 6.216127e-06, 5.2995656e-06, 4.5501676e-07, 3.6453769e-06, 5.0801686e-06, 4.867436e-07, 1.178599e-06, 4.8339925e-06, 5.132204e-07, -1.1710715e-06, 4.564241e-06, 5.3451646e-07, -3.392044e-06, 4.2741303e-06, 5.507361e-07, -5.47428e-06, 3.9668657e-06, 5.6201645e-07, -7.4092886e-06, 3.6456172e-06, 5.6852446e-07, -9.190113e-06, 3.313498e-06, 5.7045446e-07, -1.0811303e-05, 2.9735443e-06, 5.680249e-07, -1.2268877e-05, 2.628696e-06, 5.6147593e-07, -1.3560282e-05, 2.2817796e-06, 5.510661e-07, -1.4684335e-05, 1.935494e-06, 5.370697e-07, -1.5641166e-05, 1.5923952e-06, 5.1977406e-07, -1.6432148e-05, 1.2548853e-06, 4.9947624e-07, -1.7059821e-05, 9.252026e-07, 4.7648095e-07, -1.752782e-05, 6.0541254e-07, 4.510973e-07, -1.7840786e-05, 2.9740156e-07, 4.236366e-07, -1.8004284e-05, 2.872007e-09, 3.944099e-07, -1.8024713e-05, -2.7666135e-07, 3.6372558e-07, -1.7909213e-05, -5.3987293e-07, 3.3188715e-07, -1.7665578e-05, -7.856268e-07, 2.9919138e-07, -1.7302164e-05, -1.0129753e-06, 2.6592633e-07, -1.6827795e-05, -1.2211567e-06, 2.3236957e-07, -1.6251674e-05, -1.4095913e-06, 1.9878682e-07, -1.5583299e-05, -1.5778766e-06, 1.654304e-07, -1.4832369e-05, -1.7257813e-06, 1.3253809e-07, -1.4008711e-05, -1.8532382e-06, 1.00332116e-07, -1.3122193e-05, -1.9603362e-06, 6.901824e-08, -1.2182649e-05, -2.0473126e-06, 3.8785075e-08, -1.1199809e-05, -2.1145418e-06, 9.803556e-09, -1.018323e-05, -2.162528e-06, -1.7773452e-08, -9.142238e-06, -2.191893e-06, -4.3811365e-08, -8.085861e-06, -2.203366e-06, -6.819396e-08, -7.0227857e-06, -2.197773e-06, -9.082333e-08, -5.961305e-06, -2.1760256e-06, -1.1161961e-07, -4.909277e-06, -2.13911e-06, -1.3052077e-07, -3.8740886e-06, -2.088075e-06, -1.4748207e-07, -2.862625e-06, -2.0240216e-06, -1.6247554e-07, -1.8812433e-06, -1.9480922e-06, -1.754894e-07, -9.357506e-07, -1.8614601e-06, -1.8652722e-07, -3.139061e-08, -1.7653184e-06, -1.9560716e-07, 8.271681e-07, -1.6608706e-06, -2.0276114e-07, 1.6358373e-06, -1.549321e-06, -2.0803381e-07, 2.3911102e-06, -1.4318658e-06, -2.1148162e-07, 3.090058e-06, -1.3096843e-06, -2.1317179e-07, 3.7303223e-06, -1.1839309e-06, -2.1318127e-07, 4.3101036e-06, -1.0557281e-06, -2.1159562e-07, 4.8281468e-06, -9.2615954e-07, -2.08508e-07, 5.2837217e-06, -7.9626363e-07, -2.0401805e-07, 5.676604e-06, -6.670286e-07, -1.9823081e-07, 6.0070474e-06, -5.3938714e-07, -1.9125567e-07, 6.2757613e-06, -4.1421265e-07, -1.832053e-07, 6.48388e-06, -2.9231558e-07, -1.7419472e-07, 6.632934e-06, -1.7444049e-07, -1.6434025e-07, 6.7248156e-06, -6.126401e-08, -1.5375856e-07, 6.7617502e-06, 4.660685e-08, -1.4256588e-07, 6.74626e-06, 1.486357e-07, -1.3087701e-07, 6.6811303e-06, 2.4435718e-07, -1.18804664e-07, 6.5693766e-06, 3.3337676e-07, -1.0645866e-07, 6.4142087e-06, 4.1537018e-07, -9.3945275e-08, 6.218998e-06, 4.9008213e-07, -8.1366615e-08, 5.987243e-06, 5.5732494e-07, -6.882008e-08, 5.7225384e-06, 6.169762e-07, -5.639785e-08, 5.428541e-06, 6.689765e-07, -4.4186507e-08, 5.1089405e-06, 7.133268e-07, -3.226662e-08, 4.767431e-06, 7.500851e-07, -2.071248e-08, 4.407682e-06, 7.7936323e-07, -9.591865e-09, 4.033311e-06, 8.013234e-07, 1.0341494e-09, 3.647863e-06, 8.16174e-07, 1.1111295e-08, 3.254783e-06, 8.241662e-07, 2.0592173e-08, 2.857399e-06, 8.255896e-07, 2.9436261e-08, 2.4589015e-06, 8.2076815e-07, 3.760986e-08, 2.0623258e-06, 8.1005595e-07, 4.5085997e-08, 1.6705397e-06, 7.9383324e-07, 5.18443e-08, 1.2862281e-06, 7.725019e-07, 5.7870793e-08, 9.118834e-07, 7.464817e-07, 6.3157685e-08, 5.497967e-07, 7.162061e-07, 6.770313e-08, 2.0205074e-07, 6.821181e-07, 7.151089e-08, -1.2948513e-07, 6.4466695e-07, 7.4590076e-08, -4.4315803e-07, 6.0430386e-07, 7.695477e-08, -7.3753273e-07, 5.6147894e-07, 7.8623685e-08, -1.0113915e-06, 5.166379e-07, 7.961978e-08, -1.263732e-06, 4.702186e-07, 7.996989e-08, -1.4937638e-06, 4.2264858e-07, 7.9704286e-08, -1.7009036e-06, 3.743421e-07, 7.8856324e-08, -1.884769e-06, 3.2569793e-07, 7.746201e-08, -2.045171e-06, 2.770969e-07, 7.555959e-08, -2.1821056e-06, 2.2890023e-07, 7.3189184e-08, -2.2957447e-06, 1.814477e-07, 7.039234e-08, -2.3864256e-06, 1.3505617e-07, 6.7211694e-08, -2.4546398e-06, 9.001848e-08, 6.3690585e-08, -2.501022e-06, 4.6602395e-08, 5.987268e-08, -2.526338e-06, 5.0499254e-09, 5.5801646e-08, -2.5314714e-06, -3.4423177e-08, 5.1520807e-08, -2.5174122e-06, -7.162771e-08, 4.7072866e-08, -2.4852436e-06, -1.0640106e-07, 4.2499593e-08, -2.4361286e-06, -1.3860708e-07, 3.784156e-08, -2.371298e-06, -1.6813577e-07, 3.3137916e-08, -2.2920374e-06, -1.9490273e-07, 2.842615e-08, -2.1996743e-06, -2.188485e-07, 2.3741912e-08, -2.0955672e-06, -2.399378e-07, 1.9118817e-08, -1.981093e-06, -2.5815842e-07, 1.4588318e-08, -1.8576355e-06, -2.7352033e-07, 1.0179574e-08, -1.7265759e-06, -2.8605427e-07, 5.9193446e-09, -1.5892814e-06, -2.958106e-07, 1.8319178e-09, -1.4470963e-06, -3.0285787e-07, -2.0609479e-09, -1.301333e-06, -3.0728143e-07, -5.7400578e-09, -1.1532638e-06, -3.0918181e-07, -9.188792e-09, -1.0041133e-06, -3.0867344e-07, -1.23931025e-08, -8.55052e-07, -3.0588276e-07, -1.5341481e-08, -7.0718994e-07, -3.0094697e-07, -1.8024922e-08, -5.6157165e-07, -2.9401224e-07, -2.0436858e-08, -4.1917178e-07, -2.8523226e-07, -2.2573087e-08, -2.808912e-07, -2.7476668e-07, -2.4431682e-08, -1.4755398e-07, -2.6277962e-07, -2.601289e-08, -1.9905396e-08, -2.4943827e-07, -2.7319022e-08, 1.01389844e-07, -2.3491137e-07, -2.8354323e-08, 2.1574841e-07, -2.1936793e-07, -2.9124852e-08, 3.2266857e-07, -2.0297597e-07, -2.9638334e-08, 4.217297e-07, -1.859013e-07, -2.990403e-08, 5.125915e-07, -1.6830634e-07, -2.9932576e-08, 5.949922e-07, -1.5034921e-07, -2.9735835e-08, 6.687466e-07, -1.321826e-07, -2.9326761e-08, 7.3374383e-07, -1.1395306e-07, -2.871923e-08, 7.8994384e-07, -9.580006e-08, -2.7927895e-08, 8.373746e-07, -7.7855475e-08, -2.6968037e-08, 8.761282e-07, -6.0242854e-08, -2.585542e-08, 9.0635683e-07, -4.3076984e-08, -2.4606143e-08, 9.282688e-07, -2.6463466e-08, -2.3236513e-08, 9.421238e-07, -1.0498387e-08, -2.1762903e-08, 9.4822883e-07, 4.7319095e-09, -2.0201625e-08, 9.4693297e-07, 1.915097e-08, -1.8568825e-08, 9.386229e-07, 3.2692306e-08, -1.6880353e-08, 9.237181e-07, 4.5299377e-08, -1.5151672e-08, 9.02666e-07, 5.692551e-08, -1.3397756e-08, 8.759371e-07, 6.753374e-08, -1.1633006e-08, 8.440204e-07, 7.70966e-08, -9.871169e-09, 8.07419e-07, 8.559585e-08, -8.125271e-09, 7.6664503e-07, 9.302211e-08, -6.4075563e-09, 7.2221604e-07, 9.937451e-08, -4.729432e-09, 6.7465044e-07, 1.04660266e-07, -3.1014293e-09, 6.244636e-07, 1.08894184e-07, -1.5331689e-09, 5.7216437e-07, 1.120982e-07, -3.3333485e-11, 5.182514e-07, 1.1430081e-07, 1.3903477e-09, 4.6320997e-07, 1.15536565e-07, 2.7311087e-09, 4.075092e-07, 1.1584548e-07, 3.9831485e-09, 3.515991e-07, 1.15272464e-07, 5.1416245e-09, 2.9590845e-07, 1.13866726e-07, 6.2026406e-09, 2.408424e-07, 1.11681196e-07, 7.1632287e-09, 1.8678092e-07, 1.0877194e-07, 8.021321e-09};
endpackage
`endif
