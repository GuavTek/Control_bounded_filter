`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam N = 4;
	localparam real hf[0:1599] = {7.1762974e-05, -5.8527927e-05, 9.9383715e-06, -5.0584856e-07, 4.3618355e-05, -5.39981e-05, 1.0120038e-05, -6.3796455e-07, 1.7815462e-05, -4.9173424e-05, 1.0195152e-05, -7.6347726e-07, -5.5166706e-06, -4.4127435e-05, 1.0165587e-05, -8.805901e-07, -2.6285741e-05, -3.8933307e-05, 1.0034716e-05, -9.876971e-07, -4.4435714e-05, -3.366279e-05, 9.807299e-06, -1.083404e-06, -5.994587e-05, -2.8385251e-05, 9.489345e-06, -1.1665433e-06, -7.282939e-05, -2.3166793e-05, 9.087969e-06, -1.236186e-06, -8.313153e-05, -1.8069457e-05, 8.61123e-06, -1.2916474e-06, -9.092737e-05, -1.3150527e-05, 8.067965e-06, -1.332489e-06, -9.631937e-05, -8.46194e-06, 7.467616e-06, -1.3585155e-06, -9.943447e-05, -4.0498053e-06, 6.82006e-06, -1.3697687e-06, -0.000100421144, 4.5966278e-08, 6.1354367e-06, -1.3665159e-06, -9.944621e-05, 3.791922e-06, 5.4239786e-06, -1.3492376e-06, -9.6691576e-05, 7.161213e-06, 4.6958535e-06, -1.3186091e-06, -9.235089e-05, 1.013364e-05, 3.961009e-06, -1.2754826e-06, -8.662626e-05, 1.269559e-05, 3.2290359e-06, -1.2208651e-06, -7.972499e-05, 1.4839886e-05, 2.509035e-06, -1.1558957e-06, -7.185638e-05, 1.6565538e-05, 1.8095083e-06, -1.0818213e-06, -6.3228785e-05, 1.7877426e-05, 1.1382558e-06, -9.999726e-07, -5.404669e-05, 1.8785906e-05, 5.02296e-07, -9.117384e-07, -4.4508157e-05, 1.9306353e-05, -9.2201866e-08, -8.1854165e-07, -3.4802397e-05, 1.9458661e-05, -6.399665e-07, -7.21815e-07, -2.5107656e-05, 1.9266696e-05, -1.1366574e-06, -6.22978e-07, -1.5589374e-05, 1.875773e-05, -1.5788805e-06, -5.234154e-07, -6.398628e-06, 1.796184e-05, -1.96419e-06, -4.244572e-07, 2.3291238e-06, 1.691132e-05, -2.2910729e-06, -3.273605e-07, 1.0474995e-05, 1.564007e-05, -2.5589216e-06, -2.3329352e-07, 1.7937331e-05, 1.418302e-05, -2.7679928e-06, -1.4332173e-07, 2.463208e-05, 1.2575553e-05, -2.919356e-06, -5.839666e-08, 3.0492878e-05, 1.0852968e-05, -3.014832e-06, 2.065315e-08, 3.5470883e-05, 9.049966e-06, -3.0569222e-06, 9.3128584e-08, 3.9534356e-05, 7.200182e-06, -3.0487333e-06, 1.5846393e-07, 4.2668013e-05, 5.3357617e-06, -2.9938944e-06, 2.162286e-07, 4.48722e-05, 3.4869815e-06, -2.8964735e-06, 2.6612634e-07, 4.6161855e-05, 1.6819226e-06, -2.7608899e-06, 3.0799262e-07, 4.656535e-05, -5.3801653e-08, -2.5918273e-06, 3.4178964e-07, 4.6123205e-05, -1.6972667e-06, -2.3941482e-06, 3.675999e-07, 4.4886685e-05, -3.228402e-06, -2.1728106e-06, 3.8561797e-07, 4.2916356e-05, -4.630104e-06, -1.9327877e-06, 3.961409e-07, 4.028058e-05, -5.8882965e-06, -1.6789926e-06, 3.9955765e-07, 3.7053993e-05, -6.9919456e-06, -1.4162101e-06, 3.963375e-07, 3.3315995e-05, -7.933023e-06, -1.1490325e-06, 3.8701776e-07, 2.9149262e-05, -8.70643e-06, -8.818039e-07, 3.721914e-07, 2.4638312e-05, -9.309884e-06, -6.18572e-07, 3.5249414e-07, 1.9868125e-05, -9.743769e-06, -3.6304726e-07, 3.2859182e-07, 1.4922865e-05, -1.0010952e-05, -1.18570064e-07, 3.0116803e-07, 9.88468e-06, -1.0116587e-05, 1.1191387e-07, 2.709122e-07, 4.832618e-06, -1.0067884e-05, 3.2587047e-07, 2.3850833e-07, -1.5834674e-07, -9.873874e-06, 5.211867e-07, 2.0462451e-07, -5.018154e-06, -9.545153e-06, 6.961725e-07, 1.6990337e-07, -9.682383e-06, -9.093637e-06, 8.4955644e-07, 1.3495368e-07, -1.4092844e-05, -8.532291e-06, 9.804747e-07, 1.00342966e-07, -1.8198041e-05, -7.8748835e-06, 1.0884548e-06, 6.659128e-08, -2.1953509e-05, -7.1357326e-06, 1.1733943e-06, 3.4166302e-08, -2.5322028e-05, -6.3294688e-06, 1.2355349e-06, 3.4795655e-09, -2.8273727e-05, -5.470805e-06, 1.275434e-06, -2.5116062e-08, -3.078606e-05, -4.5743254e-06, 1.293933e-06, -5.132775e-08, -3.284371e-05, -3.6542897e-06, 1.2921232e-06, -7.492294e-08, -3.443836e-05, -2.7244564e-06, 1.2713111e-06, -9.572854e-08, -3.5568417e-05, -1.797924e-06, 1.2329833e-06, -1.1362918e-07, -3.6238645e-05, -8.8699625e-07, 1.17877e-06, -1.2856457e-07, -3.6459736e-05, -3.0653016e-09, 1.1104111e-06, -1.4052611e-07, -3.6247824e-05, 8.4348255e-07, 1.0297221e-06, -1.4955293e-07, -3.5623973e-05, 1.6433406e-06, 9.3856187e-07, -1.5572728e-07, -3.4613622e-05, 2.388336e-06, 8.3880326e-07, -1.5916963e-07, -3.3245997e-05, 3.0714632e-06, 7.323048e-07, -1.600335e-07, -3.1553536e-05, 3.6869014e-06, 6.2088606e-07, -1.5849997e-07, -2.9571293e-05, 4.2300135e-06, 5.0630524e-07, -1.5477247e-07, -2.7336335e-05, 4.69733e-06, 3.902399e-07, -1.4907117e-07, -2.4887193e-05, 5.086519e-06, 2.7427075e-07, -1.4162802e-07, -2.2263279e-05, 5.3963463e-06, 1.5986811e-07, -1.326816e-07, -1.9504363e-05, 5.6266185e-06, 4.838156e-08, -1.2247267e-07, -1.665006e-05, 5.7781253e-06, -5.896778e-08, -1.11239736e-07, -1.373936e-05, 5.8525693e-06, -1.6109232e-07, -9.921538e-08, -1.0810192e-05, 5.8524893e-06, -2.5704063e-07, -8.6622855e-08, -7.89902e-06, 5.7811844e-06, -3.4599788e-07, -7.367326e-08, -5.040486e-06, 5.6426297e-06, -4.2728425e-07, -6.056325e-08, -2.2670938e-06, 5.4413945e-06, -5.0035175e-07, -4.747317e-08, 3.9106783e-07, 5.1825555e-06, -5.6477955e-07, -3.4565804e-08, 2.9065584e-06, 4.871615e-06, -6.202681e-07, -2.1985565e-08, 5.2547775e-06, 4.5144193e-06, -6.666322e-07, -9.858122e-09, 7.414116e-06, 4.117076e-06, -7.03794e-07, 1.7095175e-09, 9.366067e-06, 3.6858778e-06, -7.3177443e-07, 1.262856e-08, 1.1095303e-05, 3.2272287e-06, -7.506858e-07, 2.2827649e-08, 1.2589709e-05, 2.7475728e-06, -7.60723e-07, 3.225181e-08, 1.3840387e-05, 2.2533272e-06, -7.6215593e-07, 4.0861167e-08, 1.4841629e-05, 1.7508199e-06, -7.5532125e-07, 4.8629516e-08, 1.5590856e-05, 1.2462306e-06, -7.40615e-07, 5.5542746e-08, 1.6088528e-05, 7.455371e-07, -7.184858e-07, 6.159724e-08, 1.633804e-05, 2.5446525e-07, -6.8942774e-07, 6.679825e-08, 1.6345564e-05, -2.2155695e-07, -6.5397444e-07, 7.115831e-08, 1.6119917e-05, -6.7744065e-07, -6.126935e-07, 7.469572e-08, 1.567236e-05, -1.1084736e-06, -5.661809e-07, 7.7433185e-08, 1.5016408e-05, -1.510353e-06, -5.1505646e-07, 7.939655e-08, 1.4167622e-05, -1.8792148e-06, -4.5995927e-07, 8.0613724e-08, 1.3143379e-05, -2.211659e-06, -4.015433e-07, 8.1113804e-08, 1.1962637e-05, -2.5047705e-06, -3.4047358e-07, 8.0926384e-08, 1.0645684e-05, -2.756136e-06, -2.7742223e-07, 8.008104e-08, 9.213888e-06, -2.963857e-06, -2.1306467e-07, 7.860703e-08, 7.689438e-06, -3.1265592e-06, -1.4807578e-07, 7.65332e-08, 6.0950724e-06, -3.2433963e-06, -8.312596e-08, 7.3888e-08, 4.4538265e-06, -3.3140511e-06, -1.8877099e-08, 7.0699755e-08, 2.7887604e-06, -3.338732e-06, 4.402163e-08, 6.69969e-08, 1.1227004e-06, -3.3181636e-06, 1.0493817e-07, 6.2808496e-08, -5.220158e-07, -3.253575e-06, 1.632622e-07, 5.816469e-08, -2.1237872e-06, -3.1466825e-06, 2.1840992e-07, 5.3097274e-08, -3.6619886e-06, -2.9996672e-06, 2.6982903e-07, 4.7640235e-08, -5.117195e-06, -2.8151494e-06, 3.1700384e-07, 4.1830287e-08, -6.4713963e-06, -2.5961579e-06, 3.5946036e-07, 3.5707366e-08, -7.70819e-06, -2.3460943e-06, 3.9677155e-07, 2.9315023e-08, -8.812962e-06, -2.0686946e-06, 4.285623e-07, 2.2700748e-08, -9.773036e-06, -1.7679856e-06, 4.5451435e-07, 1.591614e-08, -1.0577818e-05, -1.4482381e-06, 4.7437086e-07, 9.016965e-09, -1.1218896e-05, -1.1139174e-06, 4.879406e-07, 2.063049e-09, -1.169013e-05, -7.6962976e-07, 4.951017e-07, -4.8819833e-09, -1.1987705e-05, -4.2006778e-07, 4.9580444e-07, -1.1751135e-08, -1.2110164e-05, -6.995334e-08, 4.900738e-07, -1.847462e-08, -1.2058406e-05, 2.7602024e-07, 4.78011e-07, -2.4980592e-08, -1.18356575e-05, 6.132467e-07, 4.5979374e-07, -3.1196034e-08, -1.1447412e-05, 9.372647e-07, 4.356763e-07, -3.704776e-08, -1.0901349e-05, 1.243815e-06, 4.0598755e-07, -4.24635e-08, -1.02072145e-05, 1.5288953e-06, 3.7112872e-07, -4.7373128e-08, -9.376679e-06, 1.788813e-06, 3.3156974e-07, -5.170987e-08, -8.423173e-06, 2.0202342e-06, 2.8784427e-07, -5.5411594e-08, -7.3616966e-06, 2.2202282e-06, 2.4054415e-07, -5.8422085e-08, -6.208603e-06, 2.3863079e-06, 1.9031224e-07, -6.069226e-08, -4.981372e-06, 2.5164638e-06, 1.3783475e-07, -6.2181364e-08, -3.6983636e-06, 2.6091925e-06, 8.383251e-08, -6.285803e-08, -2.378558e-06, 2.6635182e-06, 2.905142e-08, -6.270121e-08, -1.0412887e-06, 2.6790065e-06, -2.574763e-08, -6.170105e-08, 2.9403114e-07, 2.6557716e-06, -7.979936e-08, -5.985943e-08, 1.6081818e-06, 2.594475e-06, -1.3234502e-07, -5.719046e-08, 2.88241e-06, 2.4963176e-06, -1.8264348e-07, -5.372068e-08, 4.098694e-06, 2.3630216e-06, -2.2998225e-07, -4.9489064e-08, 5.239998e-06, 2.1968071e-06, -2.7368836e-07, -4.4546805e-08, 6.290515e-06, 2.00036e-06, -3.1313866e-07, -3.8956838e-08, 7.2358903e-06, 1.7767926e-06, -3.4776977e-07, -3.279315e-08, 8.063421e-06, 1.5295994e-06, -3.770871e-07, -2.6139872e-08, 8.762236e-06, 1.2626043e-06, -4.0067295e-07, -1.909015e-08, 9.323449e-06, 9.799045e-07, -4.1819348e-07, -1.174482e-08, 9.740277e-06, 6.858095e-07, -4.2940462e-07, -4.2109125e-09, 1.00081315e-05, 3.8477646e-07, -4.3415642e-07, 3.3999863e-09, 1.0124675e-05, 8.134348e-08, -4.3239595e-07, 1.0973502e-08, 1.0089846e-05, -2.1993922e-07, -4.2416897e-07, 1.839432e-08, 9.905847e-06, -5.1457795e-07, -4.0961962e-07, 2.55481e-08, 9.577098e-06, -7.982038e-07, -3.8898875e-07, 3.2323392e-08, 9.110161e-06, -1.0666389e-06, -3.626107e-07, 3.8613557e-08, 8.513622e-06, -1.3159599e-06, -3.309084e-07, 4.4318615e-08, 7.797956e-06, -1.5425582e-06, -2.9438698e-07, 4.9347012e-08, 6.9753505e-06, -1.7431935e-06, -2.536262e-07, 5.361729e-08, 6.059512e-06, -1.915044e-06, -2.0927148e-07, 5.7059534e-08, 5.0654435e-06, -2.0557486e-06, -1.6202353e-07, 5.961672e-08, 4.009206e-06, -2.1634412e-06, -1.12627575e-07, 6.1245785e-08, 2.9076643e-06, -2.2367792e-06, -6.186136e-08, 6.1918485e-08, 1.7782195e-06, -2.2749614e-06, -1.0522686e-08, 6.162202e-08, 6.3853537e-07, -2.2777392e-06, 4.058337e-08, 6.035935e-08, -4.9373824e-07, -2.2454176e-06, 9.065748e-08, 5.8149297e-08, -1.6012411e-06, -2.1788471e-06, 1.3891898e-07, 5.5026295e-08, -2.667172e-06, -2.0794096e-06, 1.8461853e-07, 5.103992e-08, -3.6755478e-06, -1.9489908e-06, 2.2705026e-07, 4.6254137e-08, -4.611448e-06, -1.7899505e-06, 2.6556322e-07, 4.074627e-08, -5.461242e-06, -1.60508e-06, 2.9957195e-07, 3.4605755e-08, -6.2127933e-06, -1.3975562e-06, 3.2856585e-07, 2.793266e-08, -6.85564e-06, -1.1708879e-06, 3.5211747e-07, 2.0836026e-08, -7.3811448e-06, -9.2885784e-07, 3.6988928e-07, 1.3432016e-08, -7.782618e-06, -6.7545966e-07, 3.81639e-07, 5.84196e-09, -8.055404e-06, -4.1483224e-07, 3.8722322e-07, -1.8097063e-09, -8.196942e-06, -1.5119203e-07, 3.865995e-07, -9.397564e-09, -8.206782e-06, 1.11235785e-07, 3.798267e-07, -1.6797353e-08, -8.086577e-06, 3.6828575e-07, 3.6706345e-07, -2.3888104e-08, -7.840031e-06, 6.159193e-07, 3.4856532e-07, -3.05542e-08, -7.472824e-06, 8.502895e-07, 3.2467997e-07, -3.6687364e-08, -6.992499e-06, 1.0678018e-06, 2.95841e-07, -4.2188503e-08, -6.4083206e-06, 1.2651712e-06, 2.625602e-07, -4.6969397e-08, -5.7311076e-06, 1.4394727e-06, 2.2541877e-07, -5.0954203e-08, -4.973043e-06, 1.5881861e-06, 1.8505706e-07, -5.408073e-08, -4.1474595e-06, 1.7092342e-06, 1.421636e-07, -5.630147e-08, -3.2686123e-06, 1.8010123e-06, 9.746332e-08, -5.7584398e-08, -2.3514351e-06, 1.8624106e-06, 5.170514e-08, -5.7913457e-08, -1.4112907e-06, 1.8928274e-06, 5.649252e-09, -5.7288798e-08, -4.6371366e-07, 1.8921745e-06, -3.9945668e-08, -5.572671e-08, 4.7584453e-07, 1.8608732e-06, -8.433522e-08, -5.325928e-08, 1.3922686e-06, 1.7998427e-06, -1.268017e-07, -4.9933796e-08, 2.2710228e-06, 1.7104795e-06, -1.6666588e-07, -4.5811827e-08, 3.098384e-06, 1.5946291e-06, -2.0329833e-07, -4.096812e-08, 3.8616568e-06, 1.4545511e-06, -2.3612942e-07, -3.5489244e-08, 4.5493694e-06, 1.292877e-06, -2.6465858e-07, -2.9472018e-08, 5.1514508e-06, 1.1125619e-06, -2.884621e-07, -2.3021803e-08, 5.6593763e-06, 9.1683256e-07, -3.0719968e-07, -1.6250612e-08, 6.066292e-06, 7.0912984e-07, -3.2061936e-07, -9.275146e-09, 6.3671037e-06, 4.9304896e-07, -3.2856104e-07, -2.2147402e-09, 6.5585427e-06, 2.7227756e-07, -3.3095836e-07, 4.810717e-09, 6.6391926e-06, 5.0533128e-08, -3.2783885e-07, 1.1682864e-08, 6.609492e-06, -1.6850002e-07, -3.1932262e-07, 1.82869e-08, 6.471699e-06, -3.8123193e-07, -3.0561938e-07, 2.4513565e-08, 6.2298313e-06, -5.8422626e-07, -2.870239e-07, 3.0260967e-08, 5.889575e-06, -7.742562e-07, -2.639103e-07, 3.5436315e-08, 5.458166e-06, -9.48356e-07, -2.3672456e-07, 3.9957445e-08, 4.9442483e-06, -1.1038679e-06, -2.0597638e-07, 4.375417e-08, 4.357709e-06, -1.238483e-06, -1.7222969e-07, 4.676939e-08, 3.709495e-06, -1.3502755e-06, -1.3609242e-07, 4.895997e-08, 3.0114154e-06, -1.4377307e-06, -9.820563e-08, 5.0297377e-08, 2.275928e-06, -1.4997646e-06, -5.9232153e-08, 5.0768048e-08, 1.5159231e-06, -1.5357372e-06, -1.9844975e-08, 5.0373476e-08, 7.4449855e-07, -1.545457e-06, 1.9284402e-08, 4.9130055e-08, -2.5263779e-08, -1.5291782e-06, 5.7497473e-08, 4.7068646e-08, -7.805187e-07, -1.4875905e-06, 9.415989e-08, 4.4233904e-08, -1.5088709e-06, -1.4218009e-06, 1.2867204e-07, 4.0683364e-08, -2.1985784e-06, -1.3333093e-06, 1.6047899e-07, 3.6486302e-08, -2.8387412e-06, -1.2239778e-06, 1.8907943e-07, 3.1722415e-08, -3.4194727e-06, -1.0959933e-06, 2.1403368e-07, 2.6480315e-08, -3.932053e-06, -9.518253e-07, 2.3497043e-07, 2.0855891e-08, -4.369058e-06, -7.941805e-07, 2.5159233e-07, 1.495056e-08, -4.724466e-06, -6.2595234e-07, 2.636802e-07, 8.8694225e-09, -4.993738e-06, -4.5016904e-07, 2.7109562e-07, 2.7193976e-09, -5.1738716e-06, -2.6993982e-07, 2.737825e-07, -3.3926755e-09, -5.2634286e-06, -8.840012e-08, 2.7176674e-07, -9.361903e-09, -5.2625323e-06, 9.134229e-08, 2.6515488e-07, -1.5087153e-08, -5.172844e-06, 2.6626043e-07, 2.5413098e-07, -2.047278e-08, -4.9975056e-06, 4.334588e-07, 2.3895245e-07, -2.5430243e-08, -4.741066e-06, 5.902213e-07, 2.199446e-07, -2.9879562e-08, -4.4093767e-06, 7.3405505e-07, 1.9749402e-07, -3.375063e-08, -4.0094715e-06, 8.6272985e-07, 1.72041e-07, -3.6984314e-08, -3.5494277e-06, 9.743129e-07, 1.4407112e-07, -3.9533365e-08, -3.0382068e-06, 1.0671969e-06, 1.1410619e-07, -4.136309e-08, -2.4854892e-06, 1.140123e-06, 8.269461e-08, -4.2451823e-08, -1.9014931e-06, 1.1921974e-06, 5.040146e-08, -4.279112e-08, -1.2967907e-06, 1.2228998e-06, 1.7798396e-08, -4.2385746e-08, -6.8211995e-07, 1.2320877e-06, -1.4546394e-08, -4.1253426e-08, -6.8196314e-08, 1.219992e-06, -4.6078068e-08, -3.942436e-08, 5.344718e-07, 1.1872071e-06, -7.6264605e-08, -3.694052e-08, 1.1157607e-06, 1.1346748e-06, -1.04605775e-07, -3.385477e-08, 1.6661e-06, 1.0636617e-06, -1.3064138e-07, -3.022978e-08, 2.1766286e-06, 9.757327e-07, -1.5395871e-07, -2.6136778e-08, 2.6393357e-06, 8.72718e-07, -1.7419906e-07, -2.1654202e-08, 3.0471842e-06, 7.5667725e-07, -1.9106312e-07, -1.6866192e-08, 3.3942167e-06, 6.298598e-07, -2.0431538e-07, -1.1861047e-08, 3.6756387e-06, 4.946622e-07, -2.1378723e-07, -6.7295916e-09, 3.8878816e-06, 3.5358383e-07, -2.1937883e-07, -1.563543e-09, 4.0286436e-06, 2.0918192e-07, -2.2105988e-07, 3.546122e-09, 4.0969057e-06, 6.402543e-08, -2.1886898e-07, 8.510768e-09, 4.0929267e-06, -7.934979e-08, -2.1291187e-07, 1.3245636e-08, 4.018217e-06, -2.1848483e-07, -2.0335851e-07, 1.7671283e-08, 3.875489e-06, -3.5103943e-07, -1.9043907e-07, 2.1714921e-08, 3.6685842e-06, -4.7483093e-07, -1.7443887e-07, 2.5311598e-08, 3.4023924e-06, -5.8786975e-07, -1.5569249e-07, 2.8405243e-08, 3.0827414e-06, -6.883909e-07, -1.3457708e-07, 3.0949526e-08, 2.7162798e-06, -7.74881e-07, -1.1150496e-07, 3.290853e-08, 2.3103455e-06, -8.461005e-07, -8.6915826e-08, 3.425725e-08, 1.8728239e-06, -9.011004e-07, -6.12685e-08, 3.4981852e-08, 1.4119996e-06, -9.3923404e-07, -3.5032517e-08, 3.5079758e-08, 9.3640404e-07, -9.60163e-07, -8.679627e-09, 3.4559527e-08, 4.5466012e-07, -9.638574e-07, 1.7324556e-08, 3.3440525e-08, -2.4670355e-08, -9.5059073e-07, 4.252872e-08, 3.1752425e-08, -4.932364e-07, -9.2093035e-07, 6.650358e-08, 2.9534503e-08, -9.4304096e-07, -8.757212e-07, 8.8849156e-08, 2.6834808e-08, -1.3665748e-06, -8.1606623e-07, 1.0920131e-07, 2.370916e-08, -1.75694e-06, -7.433024e-07, 1.2723763e-07, 2.0220039e-08, -2.1079597e-06, -6.589725e-07, 1.4268245e-07, 1.6435358e-08, -2.4142737e-06, -5.6479405e-07, 1.5531093e-07, 1.2427183e-08, -2.6714172e-06, -4.6262582e-07, 1.6495214e-07, 8.270361e-09, -2.875883e-06, -3.544323e-07, 1.7149125e-07, 4.0411603e-09, -3.025165e-06, -2.4224676e-07, 1.7487052e-07, -1.8413011e-10, -3.1177829e-06, -1.2813402e-07, 1.7508938e-07, -4.3305537e-09, -3.1532893e-06, -1.4153112e-08, 1.7220343e-07, -8.325807e-09, -3.132257e-06, 9.767913e-08, 1.6632248e-07, -1.2101491e-08, -3.0562499e-06, 2.0542316e-07, 1.5760762e-07, -1.5594267e-08, -2.9277746e-06, 3.0724985e-07, 1.4626744e-07, -1.8746913e-08, -2.7502192e-06, 4.0147083e-07, 1.3255352e-07, -2.1509242e-08, -2.5277743e-06, 4.8656614e-07, 1.16755125e-07, -2.3838888e-08, -2.265344e-06, 5.6120797e-07, 9.919336e-08, -2.570194e-08, -1.968443e-06, 6.242807e-07, 8.02149e-08, -2.70734e-08, -1.6430885e-06, 6.748971e-07, 6.0185336e-08, -2.7937492e-08, -1.2956809e-06, 7.124094e-07, 3.948225e-08, -2.8287793e-08, -9.3288355e-07, 7.364168e-07, 1.8488265e-08, -2.8127186e-08, -5.6149736e-07, 7.467674e-07, -2.4158833e-09, -2.7467655e-08, -1.8833748e-07, 7.435567e-07, -2.2858172e-08, -2.6329916e-08, 1.7988927e-07, 7.2712083e-07, -4.248179e-08, -2.4742903e-08, 5.367024e-07, 6.980261e-07, -6.0951265e-08, -2.27431e-08, 8.7595896e-07, 6.5705433e-07, -7.79581e-08, -2.037377e-08, 1.1919574e-06, 6.0518477e-07, -9.3225836e-08, -1.7684048e-08, 1.4795305e-06, 5.435725e-07, -1.0651443e-07, -1.4727967e-08, 1.7341282e-06, 4.7352484e-07, -1.176239e-07, -1.1563396e-08, 1.9518861e-06, 3.964742e-07, -1.2639723e-07, -8.2509315e-09, 2.129682e-06, 3.1395052e-07, -1.3272233e-07, -4.852767e-09, 2.2651764e-06, 2.2755151e-07, -1.3653336e-07, -1.4315347e-09, 2.35684e-06, 1.3891268e-07, -1.3781093e-07, 1.9508277e-09, 2.4039643e-06, 4.967716e-08, -1.3658168e-07, 5.2341815e-09, 2.406658e-06, -3.853415e-08, -1.3291692e-07, 8.361243e-09, 2.3658285e-06, -1.241513e-07, -1.2693056e-07, 1.1278567e-08, 2.2831503e-06, -2.0568267e-07, -1.1877621e-07, 1.3937448e-08, 2.161018e-06, -2.817404e-07, -1.08643704e-07, 1.6294713e-08, 2.0024904e-06, -3.5106342e-07, -9.675499e-08, 1.8313413e-08, 1.8112198e-06, -4.1253782e-07, -8.335953e-08, 1.9963377e-08, 1.5913756e-06, -4.652141e-07, -6.8729264e-08, 2.1221636e-08, 1.3475578e-06, -5.0832114e-07, -5.315327e-08, 2.2072724e-08, 1.0847049e-06, -5.412768e-07, -3.6932214e-08, 2.2508816e-08, 8.079978e-07, -5.6369447e-07, -2.0372688e-08, 2.2529738e-08, 5.227611e-07, -5.753867e-07, -3.781538e-09, 2.2142837e-08, 2.3436333e-07, -5.763644e-07, 1.2539708e-08, 2.1362712e-08, -5.1881397e-08, -5.668328e-07, 2.830021e-08, 2.0210825e-08, -3.308086e-07, -5.4718396e-07, 4.3224897e-08, 1.8714989e-08, -5.974944e-07, -5.1798605e-07, 5.705917e-08, 1.6908746e-08, -8.473404e-07, -4.7996946e-07, 6.957315e-08, 1.4830663e-08, -1.0761504e-06, -4.340103e-07, 8.056537e-08, 1.2523535e-08, -1.2801992e-06, -3.8111187e-07, 8.986595e-08, 1.003354e-08, -1.4562903e-06, -3.223835e-07, 9.733905e-08, 7.4093327e-09, -1.6018042e-06, -2.5901858e-07, 1.0288474e-07, 4.7011164e-09, -1.7147344e-06, -1.9227096e-07, 1.06440126e-07, 1.9597055e-09, -1.793711e-06, -1.2343104e-07, 1.07979815e-07, -7.644136e-10, -1.8380139e-06, -5.380133e-08, 1.07515646e-07, -3.4219951e-09, -1.8475719e-06, 1.5327393e-08, 1.0509581e-07, -5.965908e-09, -1.8229517e-06, 8.269956e-08, 1.00803256e-07, -8.351958e-09, -1.7653344e-06, 1.4711702e-07, 9.475354e-08, -1.05396385e-08, -1.6764811e-06, 2.0745982e-07, 8.70921e-08, -1.2492806e-08, -1.5586897e-06, 2.627052e-07, 7.799102e-08, -1.4180257e-08, -1.4147415e-06, 3.1194438e-07, 6.76454e-08, -1.5576212e-08, -1.2478406e-06, 3.5439697e-07, 5.626936e-08, -1.6660689e-08, -1.0615468e-06, 3.8942278e-07, 4.4091735e-08, -1.7419756e-08, -8.597028e-07, 4.1653078e-07, 3.1351632e-08, -1.784569e-08, -6.463585e-07, 4.3538523e-07, 1.829386e-08, -1.793699e-08, -4.2569175e-07, 4.4580878e-07, 5.1643267e-09, -1.7698309e-08, -2.0192967e-07, 4.4778255e-07, -7.794487e-09, -1.7140243e-08, 2.0730567e-08, 4.414436e-07, -2.03479e-08, -1.6279039e-08, 2.3819804e-07, 4.2707907e-07, -3.2273192e-08, -1.5136191e-08, 4.4656144e-07, 4.0511827e-07, -4.3363475e-08, -1.3737955e-08, 6.421574e-07, 3.7612173e-07, -5.3431172e-08, -1.2114775e-08, 8.2163314e-07, 3.407686e-07, -6.2311116e-08, -1.0300659e-08, 9.82002e-07, 2.998416e-07, -6.9863155e-08, -8.332485e-09, 1.1206913e-06, 2.542107e-07, -7.5974256e-08, -6.2492744e-09, 1.2355815e-06, 2.048155e-07, -8.056008e-08, -4.0914365e-09, 1.3250365e-06, 1.5264632e-07, -8.356597e-08, -1.9000046e-09, 1.3879238e-06, 9.872514e-08, -8.496744e-08, 2.8413066e-10, 1.4236261e-06, 4.4086057e-08, -8.477002e-08, 2.420968e-09, 1.4320423e-06, -1.0244001e-08, -8.300862e-08, 4.4721147e-09, 1.4135784e-06, -6.326412e-08, -7.974629e-08, 6.401462e-09, 1.3691314e-06, -1.14017375e-07, -7.5072606e-08, 8.175808e-09, 1.3000616e-06, -1.6160764e-07, -6.910144e-08, 9.765413e-09, 1.2081595e-06, -2.0521504e-07, -6.196845e-08, 1.1144488e-08, 1.095603e-06, -2.4410954e-07, -5.3828177e-08, 1.2291592e-08, 9.649107e-07, -2.7766285e-07, -4.4850815e-08, 1.318995e-08, 8.188873e-07, -3.0535793e-07, -3.5218783e-08, 1.3827679e-08, 6.605669e-07, -3.267966e-07, -2.5123143e-08, 1.4197913e-08, 4.931518e-07, -3.417045e-07, -1.4759891e-08, 1.4298845e-08, 3.1994978e-07, -3.4993383e-07, -4.3262607e-09, 1.4133663e-08, 1.4431089e-07, -3.5146374e-07, 5.9829564e-09, 1.3710405e-08, -3.0435825e-08, -3.463982e-07, 1.597896e-08, 1.3041719e-08, -2.010437e-07, -3.3496167e-07, 2.5482326e-08, 1.2144548e-08, -3.644072e-07, -3.174928e-07, 3.4326142e-08, 1.1039741e-08, -5.176169e-07, -2.9443578e-07, 4.235887e-08, 9.751596e-09, -6.5800975e-07, -2.6633015e-07, 4.944687e-08, 8.307353e-09, -7.8321403e-07, -2.3379907e-07, 5.5476534e-08, 6.736631e-09, -8.9118777e-07, -1.9753601e-07, 6.035601e-08, 5.070844e-09, -9.802503e-07, -1.5829063e-07, 6.4016525e-08, 3.342588e-09, -1.049107e-06, -1.16853776e-07, 6.641322e-08, 1.5850151e-09, -1.0968655e-06, -7.404196e-08, 6.752553e-08, -1.6878739e-10, -1.1230451e-06, -3.0681736e-08, 6.7357114e-08, -1.8864075e-09, -1.1275773e-06, 1.2405881e-08, 6.5935374e-08, -3.5366952e-09, -1.1108002e-06, 5.4420592e-08, 6.331049e-08, -5.090316e-09, -1.0734432e-06, 9.459731e-08, 5.955403e-08, -6.520261e-09, -1.0166069e-06, 1.3221974e-07, 5.47573e-08, -7.802304e-09, -9.4173544e-07, 1.6663282e-07, 4.9029246e-08, -8.915399e-09, -8.5058247e-07, 1.9725373e-07, 4.2494104e-08, -9.842014e-09, -7.4517317e-07, 2.235815e-07, 3.528882e-08, -1.0568393e-08, -6.277611e-07, 2.452047e-07, 2.756029e-08, -1.1084739e-08, -5.0078177e-07, 2.6180754e-07, 1.9462421e-08, -1.1385329e-08, -3.6680376e-07, 2.7317395e-07, 1.1153161e-08, -1.1468543e-08, -2.2847836e-07, 2.7918972e-07, 2.7914862e-09, -1.1336824e-08, -8.84883e-08, 2.7984285e-07, -5.4655795e-09, -1.0996557e-08, 5.050293e-08, 2.752218e-07, -1.3465842e-08, -1.0457883e-08, 1.859005e-07, 2.6551197e-07, -2.1064684e-08, -9.73444e-09, 3.1522555e-07, 2.5099055e-07, -2.812762e-08, -8.843051e-09, 4.3615933e-07, 2.3201964e-07, -3.4532608e-08, -7.8033535e-09, 5.4658364e-07, 2.0903785e-07, -4.01721e-08, -6.6373866e-09, 6.4461693e-07, 1.8255078e-07, -4.4954792e-08, -5.3691362e-09, 7.2864486e-07, 1.5312035e-07, -4.8807003e-08, -4.0240593e-09, 7.973459e-07, 1.213533e-07, -5.167377e-08, -2.628581e-09, 8.497105e-07, 8.788896e-08, -5.3519493e-08, -1.2095901e-09, 8.850543e-07, 5.338678e-08, -5.432828e-08, 2.0606959e-10, 9.0302535e-07, 1.851364e-08, -5.4103875e-08, 1.5920971e-09, 9.03604e-07, -1.606879e-08, -5.2869247e-08, 2.923213e-09, 8.8709794e-07, -4.9716295e-08, -5.06658e-08, 4.175611e-09, 8.5412984e-07, -8.181384e-08, -4.7552295e-08, 5.3273737e-09, 8.0562063e-07, -1.11786576e-07, -4.3603425e-08, 6.3588477e-09, 7.4276625e-07, -1.3910983e-07, -3.8908148e-08, 7.2529667e-09, 6.670106e-07, -1.6331805e-07, -3.3567773e-08, 7.995526e-09, 5.8001416e-07, -1.8401244e-07, -2.7693849e-08, 8.575393e-09, 4.8361846e-07, -2.0086723e-07, -2.1405906e-08, 8.984662e-09, 3.7980894e-07, -2.1363446e-07, -1.4829084e-08, 9.218744e-09, 2.706746e-07, -2.2214729e-07, -8.091689e-09, 9.276395e-09, 1.5836736e-07, -2.2632156e-07, -1.3227572e-09, 9.159677e-09, 4.5060336e-08, -2.2615605e-07, 5.350375e-09, 8.873865e-09, -6.709311e-08, -2.217309e-07, 1.1804415e-08, 8.427292e-09, -1.7599952e-07, -2.1320477e-07, 1.7922344e-08, 7.831137e-09, -2.7966354e-07, -2.0081042e-07, 2.3595495e-08, 7.0991715e-09, -3.7622357e-07, -1.848491e-07, 2.8725426e-08, 6.2474568e-09, -4.6398435e-07, -1.6568364e-07, 3.322559e-08, 5.294004e-09, -5.4144596e-07, -1.4373066e-07, 3.7022733e-08, 4.2584034e-09, -6.073282e-07, -1.1945173e-07, 4.0058037e-08, 3.1614358e-09};
	localparam real hb[0:1599] = {0.00010208364, -6.269006e-05, 9.649876e-06, -3.6909174e-07, 0.00013437864, -6.6413515e-05, 9.255942e-06, -2.2979255e-07, 0.00016841153, -6.963031e-05, 8.759662e-06, -9.0155645e-08, 0.0002039128, -7.227659e-05, 8.165854e-06, 4.7539764e-08, 0.00024058236, -7.429376e-05, 7.481057e-06, 1.8097502e-07, 0.0002780923, -7.562962e-05, 6.7134974e-06, 3.0783045e-07, 0.0003160905, -7.623939e-05, 5.873025e-06, 4.25826e-07, 0.0003542044, -7.6086704e-05, 4.971017e-06, 5.327631e-07, 0.00039204565, -7.5144504e-05, 4.0202513e-06, 6.2656693e-07, 0.0004292148, -7.3395815e-05, 3.0347553e-06, 7.053278e-07, 0.00046530657, -7.083441e-05, 2.02962e-06, 7.67341e-07, 0.0004999154, -6.746529e-05, 1.0207918e-06, 8.1114433e-07, 0.0005326411, -6.3305095e-05, 2.4843066e-08, 8.3555227e-07, 0.0005630947, -5.8382215e-05, -9.4128075e-07, 8.3968644e-07, 0.0005909044, -5.273683e-05, -1.8605261e-06, 8.2300096e-07, 0.00061572145, -4.6420715e-05, -2.7160106e-06, 7.853028e-07, 0.0006372257, -3.949688e-05, -3.4913073e-06, 7.2676664e-07, 0.0006551313, -3.2038966e-05, -4.1707344e-06, 6.4794284e-07, 0.00066919165, -2.4130522e-05, -4.739638e-06, 5.497593e-07, 0.00067920424, -1.5864043e-05, -5.1846714e-06, 4.3351653e-07, 0.0006850149, -7.3398583e-06, -5.4940606e-06, 3.0087557e-07, 0.00068652106, 1.3351391e-06, -5.657849e-06, 1.5383925e-07, 0.0006836753, 1.0048923e-05, -5.668125e-06, -5.2734856e-09, 0.0006764869, 1.8685885e-05, -5.519216e-06, -1.738596e-07, 0.0006650236, 2.712849e-05, -5.207855e-06, -3.4907015e-07, 0.000649412, 3.5259018e-05, -4.733309e-06, -5.278539e-07, 0.00062983733, 4.2961365e-05, -4.097474e-06, -7.0700605e-07, 0.00060654193, 5.012286e-05, -3.3049175e-06, -8.83221e-07, 0.00057982333, 5.6636098e-05, -2.3628872e-06, -1.0531484e-06, 0.00055003114, 6.240072e-05, -1.2812701e-06, -1.2134515e-06, 0.00051756285, 6.7325156e-05, -7.250485e-08, -1.360867e-06, 0.0004828594, 7.132827e-05, 1.2485498e-06, -1.4922651e-06, 0.00044639924, 7.434085e-05, 2.6647924e-06, -1.6047088e-06, 0.00040869217, 7.6307006e-05, 4.1570997e-06, -1.6955106e-06, 0.00037027244, 7.718533e-05, 5.704586e-06, -1.762287e-06, 0.00033169106, 7.69499e-05, 7.2849016e-06, -1.8030086e-06, 0.00029350806, 7.5591066e-05, 8.874564e-06, -1.8160443e-06, 0.00025628408, 7.31159e-05, 1.0449313e-05, -1.8002007e-06, 0.00022057201, 6.954856e-05, 1.1984493e-05, -1.7547528e-06, 0.00018690834, 6.4930195e-05, 1.3455449e-05, -1.6794686e-06, 0.00015580482, 5.9318736e-05, 1.4837933e-05, -1.5746238e-06, 0.00012774018, 5.27883e-05, 1.610851e-05, -1.4410087e-06, 0.00010315213, 4.542839e-05, 1.7244964e-05, -1.2799263e-06, 8.2430095e-05, 3.734281e-05, 1.822669e-05, -1.0931789e-06, 6.590824e-05, 2.8648277e-05, 1.9035071e-05, -8.8304824e-07, 5.3859494e-05, 1.9472902e-05, 1.9653822e-05, -6.5226465e-07, 4.6490237e-05, 9.954346e-06, 2.0069307e-05, -4.039682e-07, 4.3936045e-05, 2.378515e-07, 2.0270818e-05, -1.4166177e-07, 4.6258418e-05, -9.525902e-06, 2.025081e-05, 1.3084355e-07, 5.3442633e-05, -1.9183079e-05, 2.0005085e-05, 4.094894e-07, 6.5396736e-05, -2.8579056e-05, 1.9532923e-05, 6.900366e-07, 8.195177e-05, -3.7560843e-05, 1.8837154e-05, 9.681361e-07, 0.00010286322, -4.5979534e-05, 1.7924187e-05, 1.2394029e-06, 0.0001278136, -5.36927e-05, 1.6803951e-05, 1.4994921e-06, 0.00015641634, -6.0566774e-05, 1.5489803e-05, 1.744175e-06, 0.00018822077, -6.6479275e-05, 1.3998358e-05, 1.9694146e-06, 0.00022271818, -7.1320916e-05, 1.23492755e-05, 2.1714384e-06, 0.00025934892, -7.499754e-05, 1.0564976e-05, 2.3468085e-06, 0.0002975104, -7.743181e-05, 8.67032e-06, 2.4924848e-06, 0.0003365659, -7.856469e-05, 6.6922375e-06, 2.6058838e-06, 0.0003758539, -7.835662e-05, 4.659309e-06, 2.6849293e-06, 0.00041469836, -7.67884e-05, 2.6013274e-06, 2.7280944e-06, 0.00045241867, -7.386177e-05, 5.4882224e-07, 2.7344345e-06, 0.0004883404, -6.959965e-05, -1.4674297e-06, 2.70361e-06, 0.000521806, -6.4046035e-05, -3.416904e-06, 2.6358996e-06, 0.00055218494, -5.7265574e-05, -5.2698315e-06, 2.5322001e-06, 0.0005788841, -4.934276e-05, -6.9976923e-06, 2.3940197e-06, 0.0006013573, -4.038086e-05, -8.5736965e-06, 2.2234549e-06, 0.00061911455, -3.050045e-05, -9.973237e-06, 2.0231612e-06, 0.00063172984, -1.9837744e-05, -1.1174317e-05, 1.796312e-06, 0.0006388491, -8.542574e-06, -1.215793e-05, 1.5465463e-06, 0.0006401958, 3.2238208e-06, -1.2908396e-05, 1.2779115e-06, 0.00063557667, 1.5291223e-05, -1.3413649e-05, 9.947945e-07, 0.0006248851, 2.7483036e-05, -1.3665463e-05, 7.018493e-07, 0.0006081038, 3.9619004e-05, -1.3659608e-05, 4.0391748e-07, 0.000585306, 5.1518015e-05, -1.3395958e-05, 1.05946015e-07, 0.00055665517, 6.300093e-05, -1.2878514e-05, -1.8709811e-07, 0.0005224031, 7.3893425e-05, -1.2115362e-05, -4.7031367e-07, 0.00048288712, 8.402875e-05, -1.111857e-05, -7.3895046e-07, 0.00043852543, 9.325037e-05, -9.904012e-06, -9.884924e-07, 0.0003898114, 0.00010141455, -8.4911235e-06, -1.2147368e-06, 0.00033730664, 0.0001083926, -6.9026037e-06, -1.4138684e-06, 0.00028163285, 0.000114073046, -5.164056e-06, -1.5825273e-06, 0.00022346278, 0.00011836338, -3.3035808e-06, -1.7178686e-06, 0.00016351041, 0.00012119168, -1.3513243e-06, -1.8176138e-06, 0.000102520244, 0.00012250776, 6.6100876e-07, -1.8800915e-06, 4.125627e-05, 0.00012228408, 2.7006708e-06, -1.9042687e-06, -1.9509527e-05, 0.00012051621, 4.734405e-06, -1.8897699e-06, -7.900877e-05, 0.000117223, 6.728991e-06, -1.8368854e-06, -0.00013648828, 0.00011244634, 8.651788e-06, -1.7465677e-06, -0.00019122146, 0.00010625055, 1.0471273e-05, -1.6204156e-06, -0.00024251931, 9.87214e-05, 1.2157559e-05, -1.4606484e-06, -0.0002897408, 8.9964844e-05, 1.3682887e-05, -1.2700675e-06, -0.00033230256, 8.010534e-05, 1.5022085e-05, -1.0520089e-06, -0.0003696877, 6.928392e-05, 1.615298e-05, -8.1028566e-07, -0.0004014536, 5.7656016e-05, 1.705677e-05, -5.491221e-07, -0.00042723838, 4.5389028e-05, 1.771832e-05, -2.7308087e-07, -0.00044676632, 3.265968e-05, 1.8126417e-05, 1.3016105e-08, -0.0004598519, 1.9651266e-05, 1.8273959e-05, 3.0417124e-07, -0.00046640218, 6.550787e-06, 1.815805e-05, 5.952979e-07, -0.00046641813, -6.453987e-06, 1.7780061e-05, 8.8130844e-07, -0.00045999416, -1.9177442e-05, 1.7145587e-05, 1.1572026e-06, -0.00044731636, -3.1439005e-05, 1.6264356e-05, 1.4181538e-06, -0.00042865926, -4.3065957e-05, 1.5150057e-05, 1.6595928e-06, -0.0004043812, -5.389609e-05, 1.3820111e-05, 1.8772864e-06, -0.0003749185, -6.37802e-05, 1.229537e-05, 2.06741e-06, -0.00034077838, -7.258436e-05, 1.0599765e-05, 2.2266138e-06, -0.00030253077, -8.019193e-05, 8.759908e-06, 2.3520795e-06, -0.00026079916, -8.65053e-05, 6.804643e-06, 2.4415683e-06, -0.00021625093, -9.1447284e-05, 4.7645626e-06, 2.4934584e-06, -0.00016958658, -9.4962226e-05, 2.6715036e-06, 2.5067716e-06, -0.00012152896, -9.701672e-05, 5.580146e-07, 2.481189e-06, -7.281198e-05, -9.7599936e-05, -1.5431785e-06, 2.417055e-06, -2.4169287e-05, -9.67237e-05, -3.5997116e-06, 2.3153684e-06, 2.3676963e-05, -9.442205e-05, -5.580111e-06, 2.1777655e-06, 7.002706e-05, -9.0750575e-05, -7.4543054e-06, 2.0064883e-06, 0.00011421424, -8.57853e-05, -9.194111e-06, 1.8043446e-06, 0.0001556146, -7.9621335e-05, -1.0773682e-05, 1.574658e-06, 0.00019365625, -7.237119e-05, -1.2169924e-05, 1.3212086e-06, 0.00022782743, -6.416282e-05, -1.33628455e-05, 1.048167e-06, 0.00025768383, -5.513743e-05, -1.4335877e-05, 7.6002044e-07, 0.00028285457, -4.544711e-05, -1.5076106e-05, 4.614954e-07, 0.000303047, -3.5252295e-05, -1.5574473e-05, 1.5747509e-07, 0.0003180502, -2.4719135e-05, -1.5825879e-05, -1.470847e-07, 0.00032773725, -1.4016755e-05, -1.5829246e-05, -4.4724067e-07, 0.00033206595, -3.314545e-06, -1.5587499e-05, -7.381463e-07, 0.00033107825, 7.220562e-06, -1.51074755e-05, -1.0151343e-06, 0.00032489846, 1.7426728e-05, -1.439979e-05, -1.2737951e-06, 0.00031372998, 2.7149743e-05, -1.3478617e-05, -1.5100504e-06, 0.00029785096, 3.6245394e-05, -1.2361421e-05, -1.7202212e-06, 0.00027760863, 4.4581666e-05, -1.1068643e-05, -1.9010872e-06, 0.00025341284, 5.204069e-05, -9.62333e-06, -2.0499392e-06, 0.00022572836, 5.8520473e-05, -8.050725e-06, -2.1646215e-06, 0.00019506684, 6.393629e-05, -6.377833e-06, -2.2435645e-06, 0.00016197759, 6.822185e-05, -4.6329483e-06, -2.2858073e-06, 0.00012703838, 7.133009e-05, -2.8451784e-06, -2.2910092e-06, 9.084556e-05, 7.323364e-05, -1.0439487e-06, -2.2594506e-06, 5.40042e-05, 7.392501e-05, 7.4148653e-07, -2.1920237e-06, 1.7118175e-05, 7.341638e-05, 2.4825279e-06, -2.0902107e-06, -1.921955e-05, 7.173912e-05, 4.1516973e-06, -1.9560553e-06, -5.443634e-05, 6.8943016e-05, 5.7230804e-06, -1.7921217e-06, -8.798882e-05, 6.509508e-05, 7.172737e-06, -1.6014465e-06, -0.00011937117, 6.0278275e-05, 8.4790745e-06, -1.3874828e-06, -0.0001481227, 5.4589837e-05, 9.623178e-06, -1.1540371e-06, -0.00017383453, 4.8139467e-05, 1.0589086e-05, -9.052012e-07, -0.00019615534, 4.1047333e-05, 1.1364022e-05, -6.452796e-07, -0.00021479606, 3.3441895e-05, 1.19385595e-05, -3.7871396e-07, -0.00022953349, 2.545767e-05, 1.2306737e-05, -1.1000604e-07, -0.00024021267, 1.7232887e-05, 1.2466103e-05, 1.5635973e-07, -0.00024674824, 8.907149e-06, 1.2417715e-05, 4.159924e-07, -0.00024912448, 6.1909134e-07, 1.2166061e-05, 6.646684e-07, -0.0002473943, -7.4959016e-06, 1.1718945e-05, 8.984017e-07, -0.00024167694, -1.5307889e-05, 1.1087293e-05, 1.1135089e-06, -0.00023215495, -2.269444e-05, 1.0284935e-05, 1.3066689e-06, -0.00021906976, -2.9542538e-05, 9.328321e-06, 1.4749747e-06, -0.00020271653, -3.575031e-05, 8.236202e-06, 1.6159784e-06, -0.00018343837, -4.1228504e-05, 7.0292826e-06, 1.7277273e-06, -0.0001616195, -4.5901783e-05, 5.7298375e-06, 1.8087909e-06, -0.00013767814, -4.970971e-05, 4.3613104e-06, 1.8582788e-06, -0.00011205889, -5.26075e-05, 2.947898e-06, 1.8758485e-06, -8.522467e-05, -5.4566466e-05, 1.5141285e-06, 1.8617047e-06, -5.7648675e-05, -5.5574226e-05, 8.4439684e-08, 1.8165879e-06, -2.980626e-05, -5.5634588e-05, -1.3172347e-06, 1.7417547e-06, -2.166879e-06, -5.476718e-05, -2.6678633e-06, 1.6389488e-06, 2.481366e-05, -5.3006832e-05, -3.9456936e-06, 1.5103647e-06, 5.0700583e-05, -5.0402676e-05, -5.1306024e-06, 1.358603e-06, 7.508704e-05, -4.701706e-05, -6.204409e-06, 1.1866206e-06, 9.760039e-05, -4.2924225e-05, -7.1511536e-06, 9.976739e-07, 0.00011790777, -3.820882e-05, -7.957332e-06, 7.95259e-07, 0.00013572094, -3.2964243e-05, -8.612083e-06, 5.830474e-07, 0.00015080016, -2.7290911e-05, -9.107328e-06, 3.6482007e-07, 0.00016295725, -2.1294396e-05, -9.437863e-06, 1.4440091e-07, 0.00017205777, -1.5083515e-05, -9.601392e-06, -7.441041e-08, 0.00017802206, -8.768422e-06, -9.59852e-06, -2.8790365e-07, 0.00018082549, -2.4586936e-06, -9.432686e-06, -4.925207e-07, 0.00018049768, 3.7385348e-06, -9.110056e-06, -6.8491516e-07, 0.00017712083, 9.720354e-06, -8.639367e-06, -8.6200663e-07, 0.00017082722, 1.5389756e-05, -8.031726e-06, -1.0210302e-06, 0.00016179578, 2.0657188e-05, -7.3003785e-06, -1.1595796e-06, 0.0001502481, 2.5441926e-05, -6.4604396e-06, -1.2756426e-06, 0.00013644368, 2.9673298e-05, -5.5285977e-06, -1.3676304e-06, 0.00012067457, 3.329168e-05, -4.5227953e-06, -1.4343979e-06, 0.00010325977, 3.6249305e-05, -3.4618956e-06, -1.4752565e-06, 8.453903e-05, 3.8510836e-05, -2.365339e-06, -1.4899787e-06, 6.4866595e-05, 4.0053717e-05, -1.2527929e-06, -1.4787943e-06, 4.4604745e-05, 4.086831e-05, -1.4380724e-07, -1.4423788e-06, 2.411739e-05, 4.095777e-05, 9.425242e-07, -1.3818343e-06, 3.7637064e-06, 4.033773e-05, 1.9878867e-06, -1.2986627e-06, -1.6107955e-05, 3.9035775e-05, 2.9750493e-06, -1.1947329e-06, -3.5165875e-05, 3.709069e-05, 3.888144e-06, -1.0722421e-06, -5.3100346e-05, 3.455157e-05, 4.7129165e-06, -9.336708e-07, -6.9628564e-05, 3.1476724e-05, 5.4369434e-06, -7.8173565e-07, -8.449895e-05, 2.793248e-05, 6.049815e-06, -6.193369e-07, -9.749479e-05, 2.3991834e-05, 6.543277e-06, -4.495046e-07, -0.00010843728, 1.9733054e-05, 6.9113316e-06, -2.7534313e-07, -0.00011718774, 1.5238178e-05, 7.150302e-06, -9.997521e-08, -0.00012364915, 1.0591511e-05, 7.2588464e-06, 7.3513135e-08, -0.00012776688, 5.8780874e-06, 7.2379394e-06, 2.4212636e-07, -0.00012952868, 1.1821646e-06, 7.0908054e-06, 4.0301055e-07, -0.00012896398, -3.4142374e-06, 6.822819e-06, 5.53501e-07, -0.00012614229, -7.832732e-06, 6.441367e-06, 6.911661e-07, -0.00012117121, -1.1999867e-05, 5.955677e-06, 8.138457e-07, -0.000114193535, -1.5848309e-05, 5.3766184e-06, 9.196845e-07, -0.000105383995, -1.9317902e-05, 4.7164767e-06, 1.0071594e-06, -9.49454e-05, -2.235657e-05, 3.9887086e-06, 1.0751004e-06, -8.310442e-05, -2.4921057e-05, 3.2076791e-06, 1.1227041e-06, -7.0107046e-05, -2.6977506e-05, 2.3883888e-06, 1.1495426e-06, -5.621374e-05, -2.8501843e-05, 1.5461957e-06, 1.1555627e-06, -4.16945e-05, -2.9479994e-05, 6.9653515e-07, 1.1410809e-06, -2.6823873e-05, -2.9907913e-05, -1.453556e-07, 1.1067704e-06, -1.1875931e-05, -2.979143e-05, -9.647046e-07, 1.0536426e-06, 2.880572e-06, -2.9145931e-05, -1.747458e-06, 9.830231e-07, 1.7186865e-05, -2.7995866e-05, -2.4805154e-06, 8.965221e-07, 3.0798543e-05, -2.637412e-05, -3.151944e-06, 7.959999e-07, 4.3489603e-05, -2.4321238e-05, -3.7511668e-06, 6.835297e-07, 5.505603e-05, -2.1884522e-05, -4.2691236e-06, 5.6135656e-07, 6.531896e-05, -1.9117038e-05, -4.698402e-06, 4.3185364e-07, 7.412729e-05, -1.6076552e-05, -5.033334e-06, 2.9747798e-07, 8.135971e-05, -1.28243655e-05, -5.270064e-06, 1.6072464e-07, 8.692624e-05, -9.424159e-06, -5.406577e-06, 2.4081567e-08, 9.076905e-05, -5.9407826e-06, -5.4427e-06, -1.1001481e-07, 9.2862814e-05, -2.4390733e-06, -5.3800627e-06, -2.392222e-07, 9.321437e-05, 1.0173161e-06, -5.2220344e-06, -3.6133258e-07, 9.186183e-05, 4.3670343e-06, -4.9736245e-06, -4.7430916e-07, 8.887322e-05, 7.552085e-06, -4.64136e-06, -5.763197e-07, 8.4344494e-05, 1.05188e-05, -4.2331358e-06, -6.657651e-07, 7.839719e-05, 1.3218707e-05, -3.7580426e-06, -7.4130435e-07, 7.117563e-05, 1.5609294e-05, -3.2261805e-06, -8.0187266e-07, 6.284374e-05, 1.7654644e-05, -2.6484536e-06, -8.4669597e-07, 5.358167e-05, 1.9325931e-05, -2.0363577e-06, -8.7529895e-07, 4.3582124e-05, 2.0601798e-05, -1.401759e-06, -8.8750784e-07, 3.3046566e-05, 2.1468562e-05, -7.566731e-07, -8.834475e-07, 2.2181368e-05, 2.1920303e-05, -1.1304351e-07, -8.6353367e-07, 1.1193921e-05, 2.1958793e-05, 5.174727e-07, -8.284594e-07, 2.8885455e-07, 2.1593289e-05, 1.1237101e-06, -7.791775e-07, -1.0335643e-05, 2.084021e-05, 1.6951873e-06, -7.16878e-07, -2.0491287e-05, 1.9722665e-05, 2.2222825e-06, -6.42962e-07, -3.000291e-05, 1.8269891e-05, 2.6963903e-06, -5.5901234e-07, -3.8711354e-05, 1.6516582e-05, 3.110057e-06, -4.6676126e-07, -4.6476023e-05, 1.4502136e-05, 3.4570917e-06, -3.6805616e-07, -5.3177027e-05, 1.2269826e-05, 3.7326527e-06, -2.6482385e-07, -5.8716898e-05, 9.8659275e-06, 3.933307e-06, -1.5903403e-07, -6.302187e-05, 7.3388064e-06, 4.0570653e-06, -5.2662692e-08, -6.6042696e-05, 4.737982e-06, 4.1033836e-06, 5.234378e-08, -6.7754976e-05, 2.1131987e-06, 4.0731484e-06, 1.5410346e-07, -6.815905e-05, -4.864944e-07, 3.9686265e-06, 2.508318e-07, -6.727943e-05, -3.0136262e-06, 3.7933971e-06, 3.4087208e-07, -6.516378e-05, -5.4231423e-06, 3.5522569e-06, 4.2272325e-07, -6.188154e-05, -7.673179e-06, 3.2511086e-06, 4.950639e-07, -5.752214e-05, -9.725765e-06, 2.8968293e-06, 5.56773e-07, -5.2192867e-05, -1.1547435e-05, 2.497124e-06, 6.0694634e-07, -4.6016536e-05, -1.3109745e-05, 2.0603661e-06, 6.449086e-07, -3.9128816e-05, -1.438969e-05, 1.5954323e-06, 6.702214e-07, -3.1675467e-05, -1.537001e-05, 1.111527e-06, 6.8268656e-07, -2.380939e-05, -1.603938e-05, 6.1800716e-07, 6.8234465e-07, -1.568765e-05, -1.6392498e-05, 1.2420715e-07, 6.6947e-07, -7.468458e-06, -1.6430042e-05, -3.6073234e-07, 6.44561e-07, 6.9178424e-07, -1.6158541e-05, -8.280287e-07, 6.083261e-07, 8.64135e-06, -1.5590114e-05, -1.2694117e-06, 5.6166743e-07, 1.6235905e-05, -1.4742136e-05, -1.677265e-06, 5.056598e-07, 2.3341026e-05, -1.3636799e-05, -2.0447537e-06, 4.415279e-07, 2.983449e-05, -1.2300595e-05, -2.3659338e-06, 3.7062102e-07, 3.560827e-05, -1.0763738e-05, -2.6358437e-06, 2.9438553e-07, 4.0570256e-05, -9.059519e-06, -2.8505754e-06, 2.1433664e-07, 4.46456e-05, -7.2236226e-06, -3.0073259e-06, 1.3202913e-07, 4.7777758e-05, -5.2934156e-06, -3.1044256e-06, 4.902803e-08, 4.9929135e-05, -3.3072147e-06, -3.141346e-06, -3.3120354e-08, 5.1081377e-05, -1.303552e-06, -3.1186873e-06, -1.1291652e-07, 5.1235307e-05, 6.7954437e-07, -3.0381427e-06, -1.8893442e-07, 5.041049e-05, 2.6052496e-06, -2.9024463e-06, -2.5984633e-07, 4.8644455e-05, 4.438603e-06, -2.7153003e-06, -3.244453e-07, 4.5991634e-05, 6.1471196e-06, -2.4812869e-06, -3.8166513e-07, 4.2521948e-05, 7.7013465e-06, -2.205766e-06, -4.305972e-07, 3.8319195e-05, 9.075348e-06, -1.8947596e-06, -4.7050418e-07, 3.3479173e-05, 1.0247119e-05, -1.554827e-06, -5.0083025e-07, 2.8107626e-05, 1.1198909e-05, -1.1929317e-06, -5.21208e-07, 2.2318058e-05, 1.1917476e-05, -8.16304e-07, -5.3146124e-07, 1.6229435e-05, 1.2394229e-05, -4.323018e-07, -5.3160494e-07, 9.963831e-06, 1.2625304e-05, -4.827045e-08, -5.218408e-07, 3.6440829e-06, 1.2611536e-05, 3.2859325e-07, -5.025502e-07, -2.6085488e-06, 1.23583395e-05, 6.913722e-07, -4.742837e-07, -8.67662e-06, 1.1875529e-05, 1.033552e-06, -4.3774736e-07, -1.4448637e-05, 1.1177032e-05, 1.349135e-06, -3.937868e-07, -1.982103e-05, 1.0280554e-05, 1.6327408e-06, -3.433688e-07, -2.4699943e-05, 9.207163e-06, 1.8796953e-06, -2.875612e-07, -2.90028e-05, 7.980833e-06, 2.0861034e-06, -2.2751084e-07, -3.265964e-05, 6.6279317e-06, 2.248907e-06, -1.6442118e-07, -3.5614165e-05, 5.1766783e-06, 2.365925e-06, -9.952861e-08, -3.782454e-05, 3.6565784e-06, 2.4358765e-06, -3.4078983e-08, -3.9263876e-05, 2.0978432e-06, 2.4583887e-06, 3.069569e-08, -3.992046e-05, 5.308073e-07, 2.433985e-06, 9.359987e-08, -3.9797644e-05, -1.0146432e-06, 2.3640578e-06, 1.5349598e-07, -3.8913502e-05, -2.5096238e-06, 2.250826e-06, 2.0932443e-07, -3.7300197e-05, -3.926775e-06, 2.0972777e-06, 2.6012185e-07, -3.5003075e-05, -5.2407477e-06, 1.9070992e-06, 3.0503716e-07, -3.2079573e-05, -6.42864e-06, 1.6845923e-06, 3.4334528e-07, -2.8597882e-05, -7.4703817e-06, 1.4345827e-06, 3.7445815e-07, -2.4635454e-05, -8.349056e-06, 1.1623193e-06, 3.979333e-07, -2.0277352e-05, -9.0511585e-06, 8.733677e-07, 4.1347906e-07, -1.5614502e-05, -9.566785e-06, 5.735e-07, 4.2095735e-07, -1.0741849e-05, -9.889747e-06, 2.685831e-07, 4.203833e-07, -5.756498e-06, -1.0017623e-05, -3.5533432e-08, 4.119221e-07, -7.5582375e-07, -9.9517265e-06, -3.3312648e-07, 3.9588312e-07, 4.164372e-06, -9.697011e-06, -6.1870423e-07, 3.7271144e-07, 8.911643e-06, -9.26191e-06, -8.8710493e-07, 3.4297705e-07, 1.3398584e-05, -8.658112e-06, -1.1335874e-06, 3.0736186e-07, 1.7544393e-05, -7.900278e-06, -1.3539118e-06, 2.666449e-07, 2.1276273e-05, -7.005708e-06, -1.5444105e-06, 2.2168601e-07, 2.453066e-05, -5.9939675e-06, -1.7020456e-06, 1.7340835e-07, 2.7254257e-05, -4.886475e-06, -1.8244543e-06, 1.2277991e-07, 2.9404846e-05, -3.7060634e-06, -1.9099814e-06, 7.079464e-08, 3.095189e-05, -2.476524e-06, -1.9576962e-06, 1.8453473e-08, 3.187689e-05, -1.2221394e-06, -1.9673978e-06, -3.3254565e-08, 3.217351e-05, 3.278466e-08, -1.9396045e-06, -8.3370566e-08, 3.184748e-05, 1.2643774e-06, -1.8755314e-06, -1.3098311e-07, 3.0916268e-05, 2.4496458e-06, -1.7770546e-06, -1.7524444e-07, 2.9408531e-05, 3.5668927e-06, -1.6466641e-06, -2.1538511e-07, 2.7363363e-05, 4.596103e-06, -1.4874057e-06, -2.5072697e-07, 2.4829378e-05, 5.5192904e-06, -1.3028139e-06, -2.8069417e-07, 2.1863614e-05, 6.3208013e-06, -1.0968361e-06, -3.0482204e-07, 1.8530294e-05, 6.9875673e-06, -8.737518e-07, -3.2276387e-07, 1.4899487e-05, 7.509306e-06, -6.380855e-07, -3.3429515e-07, 1.1045676e-05, 7.878665e-06, -3.9451754e-07, -3.3931556e-07, 7.046268e-06, 8.091309e-06, -1.4779337e-07, -3.3784875e-07, 2.9800765e-06, 8.145946e-06, 9.736692e-08, -3.3003948e-07, -1.0741976e-06, 8.0443015e-06, 3.3635683e-07, -3.1614894e-07, -5.0394524e-06, 7.791029e-06, 5.64768e-07, -2.965476e-07, -8.841618e-06, 7.3935717e-06, 7.784696e-07, -2.717064e-07, -1.2411007e-05, 6.8619725e-06, 9.736812e-07, -2.4218622e-07, -1.5683556e-05, 6.20864e-06, 1.1470371e-06, -2.0862564e-07, -1.8601937e-05, 5.4480724e-06, 1.2956432e-06, -1.7172769e-07, -2.1116539e-05, 4.5965458e-06, 1.4171223e-06, -1.3224556e-07, -2.3186256e-05, 3.671778e-06, 1.5096506e-06, -9.096754e-08, -2.4779132e-05, 2.692568e-06, 1.571981e-06, -4.8701708e-08, -2.5872805e-05, 1.6784231e-06, 1.6034579e-06, -6.2604064e-09, -2.6454762e-05, 6.491779e-07, 1.6040183e-06, 3.5555022e-08, -2.6522412e-05, -3.753856e-07, 1.574183e-06, 7.596906e-08, -2.6082966e-05, -1.3759102e-06, 1.5150366e-06, 1.142461e-07, -2.515313e-05, -2.3338214e-06, 1.4281976e-06, 1.497035e-07, -2.3758632e-05, -3.2316652e-06, 1.3157784e-06, 1.8172342e-07, -2.1933587e-05, -4.0534173e-06, 1.180337e-06, 2.0976339e-07, -1.9719697e-05, -4.7847625e-06, 1.0248218e-06, 2.3336499e-07, -1.7165352e-05, -5.4133347e-06, 8.525091e-07, 2.521611e-07, -1.4324592e-05, -5.928917e-06, 6.6693565e-07, 2.6588117e-07, -1.125599e-05, -6.3235993e-06, 4.7182812e-07, 2.7435456e-07, -8.021481e-06, -6.5918885e-06, 2.7102968e-07, 2.775121e-07, -4.6851233e-06, -6.73077e-06, 6.842567e-08, 2.7538556e-07, -1.311858e-06, -6.7397254e-06, -1.3213008e-07, 2.6810537e-07, 2.0337316e-06, -6.6206985e-06, -3.2688715e-07, 2.5589645e-07, 5.2886357e-06, -6.3780185e-06, -5.122673e-07, 2.3907236e-07, 8.3925825e-06, -6.018279e-06, -6.849289e-07, 2.1802799e-07, 1.1289128e-05, -5.550175e-06, -8.4182557e-07, 1.9323063e-07, 1.3926667e-05, -4.9843065e-06, -9.802585e-07, 1.6521012e-07, 1.6259315e-05, -4.3329446e-06, -1.0979217e-06, 1.3454775e-07, 1.8247698e-05, -3.6097745e-06, -1.1929379e-06, 1.0186454e-07, 1.9859572e-05, -2.829613e-06, -1.263888e-06, 6.780895e-08, 2.1070327e-05, -2.0081134e-06, -1.3098283e-06, 3.30442e-08, 2.1863327e-05, -1.1614534e-06, -1.3303022e-06, -1.7643523e-09, 2.223009e-05, -3.060251e-07, -1.3253392e-06, -3.5961733e-08, 2.2170316e-05, 5.418789e-07, -1.2954471e-06, -6.891546e-08, 2.1691769e-05, 1.36637e-06, -1.2415941e-06, -1.0002699e-07, 2.080999e-05, 2.1522567e-06, -1.1651832e-06, -1.2874239e-07, 1.9547888e-05, 2.8853178e-06, -1.068019e-06, -1.5456192e-07, 1.7935185e-05, 3.5525557e-06, -9.522662e-07, -1.7704856e-07, 1.6007747e-05, 4.142421e-06, -8.2040407e-07, -1.9583507e-07, 1.3806819e-05, 4.6450045e-06, -6.7517425e-07, -2.1062976e-07, 1.1378147e-05, 5.0522e-06, -5.1952486e-07, -2.2122063e-07, 8.7710605e-06, 5.3578256e-06, -3.5655214e-07, -2.274781e-07, 6.037475e-06, 5.557709e-06, -1.894396e-07, -2.2935593e-07, 3.2308817e-06, 5.649735e-06, -2.1397017e-08, -2.2689086e-07, 4.0531154e-07, 5.6338513e-06, 1.4440032e-07, -2.2020043e-07, -2.385688e-06, 5.512036e-06, 3.0487055e-07, -2.0947948e-07, -5.090054e-06, 5.2882287e-06, 4.5708157e-07, -1.9499517e-07, -7.658161e-06, 4.9682258e-06, 5.9830364e-07, -1.7708086e-07, -1.004372e-05, 4.55954e-06, 7.260573e-07, -1.5612873e-07, -1.2204593e-05, 4.0712334e-06, 8.3815564e-07, -1.3258145e-07, -1.4103522e-05, 3.5137218e-06, 9.327408e-07, -1.0692307e-07, -1.5708747e-05, 2.898559e-06, 1.0083135e-06, -7.96693e-08, -1.6994527e-05, 2.2381996e-06, 1.0637549e-06, -5.135729e-08, -1.7941518e-05, 1.5457531e-06, 1.0983422e-06, -2.2535275e-08, -1.8537045e-05, 8.347259e-07, 1.1117552e-06, 6.247923e-09, -1.8775228e-05, 1.1876252e-07, 1.1040759e-06, 3.4453144e-08, -1.8656996e-05, -5.8861286e-07, 1.0757806e-06, 6.156083e-08, -1.8189954e-05, -1.2742483e-06, 1.0277249e-06, 8.7080444e-08, -1.7388138e-05, -1.925605e-06, 9.611209e-07, 1.1055915e-07, -1.6271657e-05, -2.530982e-06, 8.775095e-07, 1.3158969e-07, -1.4866216e-05, -3.079724e-06, 7.787257e-07, 1.4981723e-07, -1.3202548e-05, -3.562402e-06, 6.668599e-07, 1.6494522e-07, -1.131576e-05, -3.970974e-06, 5.442145e-07, 1.767399e-07, -9.244607e-06, -4.298911e-06, 4.1325742e-07, 1.8503371e-07, -7.0307083e-06, -4.5412976e-06, 2.7657325e-07, 1.8972733e-07, -4.717722e-06, -4.6948976e-06, 1.3681297e-07, 1.9079043e-07, -2.350497e-06, -4.7581884e-06, -3.3566518e-09, 1.8826113e-07, 2.5785566e-08, -4.731364e-06, -1.413033e-07, 1.8224415e-07, 2.3664659e-06, -4.6163022e-06, -2.7447777e-07, 1.7290782e-07, 4.628232e-06, -4.416505e-06, -4.004604e-07, 1.6047983e-07, 6.769912e-06, -4.1370067e-06, -5.1700425e-07, 1.452421e-07, 8.753209e-06, -3.784256e-06, -6.2207437e-07, 1.2752456e-07, 1.0543376e-05, -3.3659733e-06, -7.138825e-07, 1.0769825e-07, 1.2109812e-05, -2.8909863e-06, -7.9091683e-07, 8.61677e-08};
endpackage
`endif
