`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam N = 5;
	localparam M = 5;
	localparam COEFF_BIAS = 48;
	localparam logic signed[63:0] Lfr[0:4] = {64'd274543124250420, 64'd274543124250420, 64'd268151763923252, 64'd268151763923252, 64'd265872740036770};
	localparam logic signed[63:0] Lfi[0:4] = {64'd34346692233416, - 64'd34346692233416, 64'd20195329106117, - 64'd20195329106117, 64'd0};
	localparam logic signed[63:0] Lbr[0:4] = {64'd274543124250420, 64'd274543124250420, 64'd268151763923252, 64'd268151763923252, 64'd265872740036770};
	localparam logic signed[63:0] Lbi[0:4] = {64'd34346692233416, - 64'd34346692233416, 64'd20195329106117, - 64'd20195329106117, 64'd0};
	localparam logic signed[63:0] Wfr[0:4] = {- 64'd6335044276, - 64'd6335044276, - 64'd8643346889, - 64'd8643346889, - 64'd11515156126};
	localparam logic signed[63:0] Wfi[0:4] = {- 64'd20839617857, 64'd20839617857, 64'd9960918574, - 64'd9960918574, 64'd0};
	localparam logic signed[63:0] Wbr[0:4] = {64'd6335044276, 64'd6335044276, 64'd8643346889, 64'd8643346889, 64'd11515156126};
	localparam logic signed[63:0] Wbi[0:4] = {64'd20839617857, - 64'd20839617857, - 64'd9960918574, 64'd9960918574, 64'd0};
	localparam logic signed[63:0] Ffr[0:4][0:99] = '{
		'{64'd12121701392631576, - 64'd5511085814118572, - 64'd179182817565032, 64'd185632095569354, - 64'd16375895597195, 64'd9325598198400832, - 64'd5657779628121171, - 64'd40473921396927, 64'd177081116710846, - 64'd19110861806506, 64'd6479371739918228, - 64'd5711846607152701, 64'd94179714416863, 64'd166074689400989, - 64'd21457354306236, 64'd3628820118258496, - 64'd5675575756494004, 64'd222828347759746, 64'd152866262543536, - 64'd23392124950551, 64'd818262431874540, - 64'd5552578715388690, 64'd343681110330425, 64'd137734852169609, - 64'd24899090569803, - 64'd1910098079483638, - 64'd5347689141144777, 64'd455128396357463, 64'd120979854632028, - 64'd25969340329378, - 64'd4516756604170016, - 64'd5066846552975130, 64'd555760686623897, 64'd102915719072728, - 64'd26601031695251, - 64'd6965427846254730, - 64'd4716966960170498, 64'd644383636433401, 64'd83866566471041, - 64'd26799180378749, - 64'd9223499631869116, - 64'd4305802725520964, 64'd720029319829657, 64'd64160840461159, - 64'd26575351094600, - 64'd11262414283044492, - 64'd3841794198979132, 64'd781963585579850, 64'd44126071739022, - 64'd25947257272679, - 64'd13057974287534080, - 64'd3333915698514529, 64'd829689542188433, 64'd24083833356644, - 64'd24938278999926, - 64'd14590570083431264, - 64'd2791518415715291, 64'd862947248610265, 64'd4344958634419, - 64'd23576909422927, - 64'd15845329057963682, - 64'd2224172784336629, 64'd881709743541835, - 64'd14794913069079, - 64'd21896140604860, - 64'd16812186111136374, - 64'd1641512772634777, 64'd886175598422222, - 64'd33059404773208, - 64'd19932800397630, - 64'd17485877338516620, - 64'd1053084447441928, 64'd876758226895624, - 64'd50195034455864, - 64'd17726852258869, - 64'd17865859526355222, - 64'd468201012480347, 64'd854072225893131, - 64'd65974370219586, - 64'd15320670114924, - 64'd17956159210960408, 64'd104193651263810, 64'd818917060201813, - 64'd80198675265970, - 64'd12758300349201, - 64'd17765156019080896, 64'd655651115491204, 64'd772258433027506, - 64'd92700018913746, - 64'd10084722786950, - 64'd17305305865232496, 64'd1178332599016474, 64'd715207709354171, - 64'd103342838972494, - 64'd7345122162380, - 64'd16592810325669880, 64'd1665109859989971, 64'd648999776694870, - 64'd112024949781757, - 64'd4584181003857},
		'{64'd12121701392629594, - 64'd5511085814118876, - 64'd179182817564926, 64'd185632095569345, - 64'd16375895597196, 64'd9325598198398734, - 64'd5657779628121486, - 64'd40473921396816, 64'd177081116710836, - 64'd19110861806506, 64'd6479371739916055, - 64'd5711846607153022, 64'd94179714416977, 64'd166074689400979, - 64'd21457354306236, 64'd3628820118256281, - 64'd5675575756494324, 64'd222828347759860, 64'd152866262543527, - 64'd23392124950551, 64'd818262431872320, - 64'd5552578715389005, 64'd343681110330538, 64'd137734852169599, - 64'd24899090569804, - 64'd1910098079485828, - 64'd5347689141145084, 64'd455128396357574, 64'd120979854632019, - 64'd25969340329379, - 64'd4516756604172144, - 64'd5066846552975423, 64'd555760686624003, 64'd102915719072719, - 64'd26601031695252, - 64'd6965427846256764, - 64'd4716966960170772, 64'd644383636433501, 64'd83866566471033, - 64'd26799180378749, - 64'd9223499631871028, - 64'd4305802725521218, 64'd720029319829750, 64'd64160840461152, - 64'd26575351094601, - 64'd11262414283046258, - 64'd3841794198979361, 64'd781963585579935, 64'd44126071739016, - 64'd25947257272679, - 64'd13057974287535680, - 64'd3333915698514730, 64'd829689542188508, 64'd24083833356638, - 64'd24938278999926, - 64'd14590570083432674, - 64'd2791518415715463, 64'd862947248610330, 64'd4344958634414, - 64'd23576909422928, - 64'd15845329057964888, - 64'd2224172784336770, 64'd881709743541889, - 64'd14794913069083, - 64'd21896140604860, - 64'd16812186111137364, - 64'd1641512772634885, 64'd886175598422265, - 64'd33059404773211, - 64'd19932800397630, - 64'd17485877338517386, - 64'd1053084447442003, 64'd876758226895655, - 64'd50195034455866, - 64'd17726852258869, - 64'd17865859526355762, - 64'd468201012480389, 64'd854072225893150, - 64'd65974370219587, - 64'd15320670114924, - 64'd17956159210960716, 64'd104193651263801, 64'd818917060201820, - 64'd80198675265970, - 64'd12758300349202, - 64'd17765156019080980, 64'd655651115491226, 64'd772258433027502, - 64'd92700018913746, - 64'd10084722786950, - 64'd17305305865232360, 64'd1178332599016527, 64'd715207709354156, - 64'd103342838972492, - 64'd7345122162380, - 64'd16592810325669532, 64'd1665109859990052, 64'd648999776694844, - 64'd112024949781754, - 64'd4584181003857},
		'{- 64'd54230251112480224, 64'd10162912064129204, - 64'd1107410074232320, 64'd66607254859419, 64'd34180873857108, - 64'd49176792574385560, 64'd10039753153409532, - 64'd1154689346203892, 64'd90659314527461, 64'd27733084614410, - 64'd44201062489677208, 64'd9853166970426098, - 64'd1189310977363184, 64'd111942322359692, 64'd21643151376508, - 64'd39333038862206016, 64'd9610067924103708, - 64'd1212123917937735, 64'd130540713330342, 64'd15924834974848, - 64'd34599287485460208, 64'd9317184474204714, - 64'd1223990268590974, 64'd146551387709459, 64'd10587949604627, - 64'd30023063481010368, 64'd8981025649058081, - 64'd1225777763232035, 64'd160081907180583, 64'd5638634772698, - 64'd25624428434944856, 64'd8607852106801811, - 64'd1218352866297295, 64'd171248769629750, 64'd1079630659773, - 64'd21420380905485056, 64'd8203651557393658, - 64'd1202574481872452, 64'd180175768485818, - 64'd3089445435503, - 64'd17424998170533344, 64'd7774118346376153, - 64'd1179288267733101, 64'd186992441354221, - 64'd6871823707512, - 64'd13649587186875850, 64'd7324636988003550, - 64'd1149321543516658, 64'd191832611612620, - 64'd10273309452191, - 64'd10102842841729462, 64'd6860269424696720, - 64'd1113478778790348, 64'd194833025629963, - 64'd13302015424023, - 64'd6791011690960054, 64'd6385745781726976, - 64'd1072537643737978, 64'd196132087331631, - 64'd15968100504470, - 64'd3718059495358866, 64'd5905458380376236, - 64'd1027245602539384, 64'd195868690963791, - 64'd18283516061774, - 64'd885840985683144, 64'd5423458769409848, - 64'd978317027246011, 64'd194181152110122, - 64'd20261761204803, 64'd1705729592333484, 64'd4943457533359528, - 64'd926430808047790, 64'd191206236283473, - 64'd21917647962927, 64'd4058508481108936, 64'd4468826636676080, - 64'd872228434262854, 64'd187078283753276, - 64'd23267077260512, 64'd6175954170621278, 64'd4002604065104876, - 64'd816312519144131, 64'd181928428675371, - 64'd24326826399042, 64'd8062962003819387, 64'd3547500529493366, - 64'd759245740666098, 64'd175883910062924, - 64'd25114348612645, 64'd9725702601620356, 64'd3105908002494394, - 64'd701550169811212, 64'd169067471673386, - 64'd25647585124212, 64'd11171464967884652, 64'd2679909865120778, - 64'd643706957498268, 64'd161596847484811, - 64'd25944789999639},
		'{- 64'd54230251112476992, 64'd10162912064129726, - 64'd1107410074232505, 64'd66607254859435, 64'd34180873857108, - 64'd49176792574382072, 64'd10039753153410084, - 64'd1154689346204088, 64'd90659314527478, 64'd27733084614411, - 64'd44201062489673520, 64'd9853166970426672, - 64'd1189310977363388, 64'd111942322359710, 64'd21643151376509, - 64'd39333038862202176, 64'd9610067924104296, - 64'd1212123917937946, 64'd130540713330360, 64'd15924834974849, - 64'd34599287485456248, 64'd9317184474205316, - 64'd1223990268591190, 64'd146551387709477, 64'd10587949604628, - 64'd30023063481006344, 64'd8981025649058686, - 64'd1225777763232252, 64'd160081907180602, 64'd5638634772698, - 64'd25624428434940792, 64'd8607852106802416, - 64'd1218352866297513, 64'd171248769629768, 64'd1079630659774, - 64'd21420380905480984, 64'd8203651557394260, - 64'd1202574481872669, 64'd180175768485837, - 64'd3089445435502, - 64'd17424998170529294, 64'd7774118346376746, - 64'd1179288267733315, 64'd186992441354239, - 64'd6871823707511, - 64'd13649587186871850, 64'd7324636988004131, - 64'd1149321543516868, 64'd191832611612637, - 64'd10273309452190, - 64'd10102842841725546, 64'd6860269424697284, - 64'd1113478778790553, 64'd194833025629980, - 64'd13302015424022, - 64'd6791011690956236, 64'd6385745781727524, - 64'd1072537643738176, 64'd196132087331647, - 64'd15968100504469, - 64'd3718059495355164, 64'd5905458380376764, - 64'd1027245602539575, 64'd195868690963806, - 64'd18283516061773, - 64'd885840985679580, 64'd5423458769410352, - 64'd978317027246194, 64'd194181152110136, - 64'd20261761204802, 64'd1705729592336900, 64'd4943457533360008, - 64'd926430808047964, 64'd191206236283487, - 64'd21917647962926, 64'd4058508481112190, 64'd4468826636676534, - 64'd872228434263020, 64'd187078283753289, - 64'd23267077260512, 64'd6175954170624356, 64'd4002604065105303, - 64'd816312519144286, 64'd181928428675384, - 64'd24326826399041, 64'd8062962003822286, 64'd3547500529493765, - 64'd759245740666244, 64'd175883910062935, - 64'd25114348612645, 64'd9725702601623068, 64'd3105908002494765, - 64'd701550169811348, 64'd169067471673397, - 64'd25647585124212, 64'd11171464967887176, 64'd2679909865121120, - 64'd643706957498394, 64'd161596847484821, - 64'd25944789999638},
		'{- 64'd83657983348648656, 64'd9541301882050548, - 64'd2521758375897227, 64'd450532855767046, - 64'd96732342708448, - 64'd79020797936577888, 64'd9012424850491996, - 64'd2381976603908496, 64'd425559693579826, - 64'd91370441900803, - 64'd74640653008692656, 64'd8512863620693828, - 64'd2249942974631240, 64'd401970800756419, - 64'd86305752754388, - 64'd70503300739072888, 64'd8040993209566270, - 64'd2125228006348184, 64'd379689446858875, - 64'd81521800743706, - 64'd66595283062773640, 64'd7595278707286637, - 64'd2007426023633749, 64'd358643154638879, - 64'd77003024530813, - 64'd62903887899153488, 64'd7174270284512957, - 64'd1896153837764640, 64'd338763464282259, - 64'd72734725347082, - 64'd59417107801755872, 64'd6776598476349133, - 64'd1791049500275656, 64'd319985710721485, - 64'd68703019180740, - 64'd56123600900239240, 64'd6400969727721226, - 64'd1691771125606240, 64'd302248813291806, - 64'd64894791614670, - 64'd53012654007306816, 64'd6046162185674793, - 64'd1597995779008066, 64'd285495077046799, - 64'd61297655167563, - 64'd50074147770629656, 64'd5711021724906348, - 64'd1509418426096217, 64'd269670005087055, - 64'd57899908999662, - 64'd47298523756408296, 64'd5394458193600728, - 64'd1425750940627034, 64'd254722121291540, - 64'd54690500852032, - 64'd44676753357501808, 64'd5095441867362750, - 64'd1346721167275121, 64'd240602802875004, - 64'd51658991095540, - 64'd42200308424987944, 64'd4813000099708417, - 64'd1272072036360875, 64'd227266122226780, - 64'd48795518772615, - 64'd39861133527624104, 64'd4546214158220341, - 64'd1201560727648924, 64'd214668697516507, - 64'd46090769521324, - 64'd37651619748974200, 64'd4294216236075956, - 64'd1134957880497448, 64'd202769551580809, - 64'd43535945277418, - 64'd35564579936968036, 64'd4056186629227557, - 64'd1072046847789146, 64'd191529978631937, - 64'd41122735655812, - 64'd33593225325384552, 64'd3831351070052028, - 64'd1012622991217009, 64'd180913418354781, - 64'd38843290918388, - 64'd31731143451212820, 64'd3618978208797132, - 64'd956493015632619, 64'd170885336982721, - 64'd36690196440209, - 64'd29972277296059848, 64'd3418377234631920, - 64'd903474340291686, 64'd161413114965480, - 64'd34656448591071, - 64'd28310905583756036, 64'd3228895628562988, - 64'd853394504951638, 64'd152465940863573, - 64'd32735431953950}};
	localparam logic signed[63:0] Ffi[0:4][0:99] = '{
		'{64'd20467974938558076, 64'd2314420005831342, - 64'd1100572195040407, 64'd32611940301810, 64'd25718338064436, 64'd21443050477604384, 64'd1584938512519100, - 64'd1095333125455362, 64'd54460373751978, 64'd23086723774012, 64'd22052921347871056, 64'd855521716972296, - 64'd1073297268587196, 64'd74727323968669, 64'd20186186535086, 64'd22300465164129556, 64'd137470719399253, - 64'd1035373115959941, 64'd93152114409092, 64'd17070752184426, 64'd22194077140263000, - 64'd558471004406560, - 64'd982684701039992, 64'd109511415021970, 64'd13795952901513, 64'd21747353734214364, - 64'd1222265263551204, - 64'd916546904696429, 64'd123621442321922, 64'd10417915813221, 64'd20978706372071724, - 64'd1844710898556169, - 64'd838438636851291, 64'd135339472368277, 64'd6992473145366, 64'd19910913597499592, - 64'd2417558109532762, - 64'd749974381600231, 64'd144564666397293, 64'd3574306983146, 64'd18570620665159952, - 64'd2933604182346382, - 64'd652874601994840, 64'd151238219516567, 64'd216140725251, 64'd16987796106745588, - 64'd3386769757322648, - 64'd548935501598846, 64'd155342853009109, - 64'd3032011815140, 64'd15195155143353004, - 64'd3772155115444260, - 64'd439998633116790, 64'd156901680272569, - 64'd6123529972295, 64'd13227559998370616, - 64'd4086076284367489, - 64'd327920830212376, 64'd155976485111869, - 64'd9015794133221, 64'd11121407183611766, - 64'd4326081085978768, - 64'd214544917552954, 64'd152665458902827, - 64'd11670711119996, 64'd8914011693259571, - 64'd4490945553935468, - 64'd101671626696035, 64'd147100449959589, - 64'd14055151693393, 64'd6642997752742528, - 64'd4580651439364955, 64'd8966887687547, 64'd139443784197307, - 64'd16141296364669, 64'd4345705342420399, - 64'd4596345791716492, 64'd115731574875758, 64'd129884720830122, - 64'd17906887251978, 64'd2058621160268606, - 64'd4540283846211505, 64'd217098744416944, 64'd118635610348398, - 64'd19335385250248, - 64'd183157983446269, - 64'd4415756666453720, 64'd311679783473965, 64'd105927824362754, - 64'd20416033275353, - 64'd2346422118907068, - 64'd4227005178100108, 64'd398238115353751, 64'd92007528088579, - 64'd21143827773211, - 64'd4400299054528418, - 64'd3979122385158311, 64'd475703229557823, 64'd77131366294058, - 64'd21519402032049},
		'{- 64'd20467974938559408, - 64'd2314420005831492, 64'd1100572195040465, - 64'd32611940301814, - 64'd25718338064436, - 64'd21443050477605440, - 64'd1584938512519208, 64'd1095333125455406, - 64'd54460373751981, - 64'd23086723774012, - 64'd22052921347871832, - 64'd855521716972364, 64'd1073297268587226, - 64'd74727323968671, - 64'd20186186535086, - 64'd22300465164130044, - 64'd137470719399280, 64'd1035373115959956, - 64'd93152114409093, - 64'd17070752184426, - 64'd22194077140263208, 64'd558471004406573, 64'd982684701039992, - 64'd109511415021970, - 64'd13795952901513, - 64'd21747353734214296, 64'd1222265263551256, 64'd916546904696416, - 64'd123621442321920, - 64'd10417915813221, - 64'd20978706372071392, 64'd1844710898556257, 64'd838438636851265, - 64'd135339472368274, - 64'd6992473145365, - 64'd19910913597499008, 64'd2417558109532883, 64'd749974381600192, - 64'd144564666397289, - 64'd3574306983146, - 64'd18570620665159136, 64'd2933604182346534, 64'd652874601994790, - 64'd151238219516562, - 64'd216140725251, - 64'd16987796106744554, 64'd3386769757322827, 64'd548935501598786, - 64'd155342853009103, 64'd3032011815141, - 64'd15195155143351782, 64'd3772155115444463, 64'd439998633116720, - 64'd156901680272563, 64'd6123529972296, - 64'd13227559998369228, 64'd4086076284367710, 64'd327920830212300, - 64'd155976485111862, 64'd9015794133222, - 64'd11121407183610242, 64'd4326081085979006, 64'd214544917552871, - 64'd152665458902820, 64'd11670711119996, - 64'd8914011693257937, 64'd4490945553935717, 64'd101671626695948, - 64'd147100449959581, 64'd14055151693393, - 64'd6642997752740813, 64'd4580651439365210, - 64'd8966887687638, - 64'd139443784197299, 64'd16141296364670, - 64'd4345705342418633, 64'd4596345791716750, - 64'd115731574875850, - 64'd129884720830115, 64'd17906887251979, - 64'd2058621160266819, 64'd4540283846211762, - 64'd217098744417036, - 64'd118635610348390, 64'd19335385250248, 64'd183157983448051, 64'd4415756666453972, - 64'd311679783474056, - 64'd105927824362747, 64'd20416033275354, 64'd2346422118908817, 64'd4227005178100352, - 64'd398238115353839, - 64'd92007528088572, 64'd21143827773212, 64'd4400299054530106, 64'd3979122385158542, - 64'd475703229557907, - 64'd77131366294051, 64'd21519402032050},
		'{- 64'd34656575565312940, - 64'd4988108285545681, 64'd1389538734008945, - 64'd379170625264187, 64'd67317163494705, - 64'd36907080549404824, - 64'd4022832490582728, 64'd1244312214721891, - 64'd356444177497412, 64'd66583219400563, - 64'd38688484455219192, - 64'd3112083068544692, 64'd1102567579945230, - 64'd333067760901026, 64'd65421398079712, - 64'd40028568385265104, - 64'd2257829886078850, 64'd965048182911008, - 64'd309270815359571, 64'd63877628016734, - 64'd40955949332034712, - 64'd1461453472484437, 64'd832401280626865, - 64'd285265862491704, 64'd61996651052703, - 64'd41499795792327800, - 64'd723786256669338, 64'd705181638932075, - 64'd261248412089143, 64'd59821795389116, - 64'd41689564127765800, - 64'd45154254508206, 64'd583855506258482, - 64'd237397002409543, 64'd57394778848132, - 64'd41554755808632264, 64'd574581140706096, 64'd468804894556953, - 64'd213873362342983, 64'd54755541201951, - 64'd41124695511916016, 64'd1135981582474870, 64'd360332108951655, - 64'd190822683616961, 64'd51942104273018, - 64'd40428329892898456, 64'd1639990698407458, 64'd258664470947135, - 64'd168373991424715, 64'd48990458414845, - 64'd39494046712652536, 64'd2087893780182719, 64'd163959183398814, - 64'd146640602148313, 64'd45934473909715, - 64'd38349513881148224, 64'd2481278467416686, 64'd76308288930206, - 64'd125720657193185, 64'd42805835763154, - 64'd37021537866946880, 64'd2821996629167747, - 64'd4256322993214, - 64'd105697722347071, 64'd39634000334883, - 64'd35535940829298876, 64'd3112127620180786, - 64'd77757901573789, - 64'd86641442516250, 64'd36446172220825, - 64'd33917455746356300, 64'd3353943063357565, - 64'd144269850470854, - 64'd68608242168432, 64'd33267299789458, - 64'd32189638743641944, 64'd3549873285442806, - 64'd203910808051241, - 64'd51642062318009, 64'd30120087777389, - 64'd30374797769297368, 64'd3702475509617544, - 64'd256839822823478, - 64'd35775125419248, 64'd27025025362152, - 64'd28493936716348648, 64'd3814403886660708, - 64'd303251651393346, - 64'd21028720080413, 64'd24000428154009, - 64'd26566714056631972, 64'd3888381425628816, - 64'd343372202987290, - 64'd7413998071185, 64'd21062492581666, - 64'd24611415025441952, 64'd3927173865649788, - 64'd377454151408487, 64'd5067223338071, 64'd18225361188348},
		'{64'd34656575565318544, 64'd4988108285546430, - 64'd1389538734009220, 64'd379170625264209, - 64'd67317163494703, 64'd36907080549409936, 64'd4022832490583405, - 64'd1244312214722141, 64'd356444177497432, - 64'd66583219400562, 64'd38688484455223808, 64'd3112083068545297, - 64'd1102567579945454, 64'd333067760901043, - 64'd65421398079711, 64'd40028568385269240, 64'd2257829886079385, - 64'd965048182911207, 64'd309270815359586, - 64'd63877628016733, 64'd40955949332038376, 64'd1461453472484904, - 64'd832401280627039, 64'd285265862491717, - 64'd61996651052702, 64'd41499795792331008, 64'd723786256669740, - 64'd705181638932225, 64'd261248412089155, - 64'd59821795389115, 64'd41689564127768560, 64'd45154254508545, - 64'd583855506258609, 64'd237397002409552, - 64'd57394778848131, 64'd41554755808634608, - 64'd574581140705816, - 64'd468804894557059, 64'd213873362342991, - 64'd54755541201951, 64'd41124695511917952, - 64'd1135981582474646, - 64'd360332108951740, 64'd190822683616967, - 64'd51942104273017, 64'd40428329892900008, - 64'd1639990698407288, - 64'd258664470947200, 64'd168373991424719, - 64'd48990458414844, 64'd39494046712653728, - 64'd2087893780182598, - 64'd163959183398862, 64'd146640602148316, - 64'd45934473909715, 64'd38349513881149088, - 64'd2481278467416612, - 64'd76308288930236, 64'd125720657193187, - 64'd42805835763154, 64'd37021537866947424, - 64'd2821996629167714, 64'd4256322993199, 64'd105697722347071, - 64'd39634000334883, 64'd35535940829299128, - 64'd3112127620180794, 64'd77757901573789, 64'd86641442516249, - 64'd36446172220825, 64'd33917455746356280, - 64'd3353943063357609, 64'd144269850470866, 64'd68608242168430, - 64'd33267299789458, 64'd32189638743641684, - 64'd3549873285442882, 64'd203910808051266, 64'd51642062318007, - 64'd30120087777389, 64'd30374797769296888, - 64'd3702475509617648, 64'd256839822823513, 64'd35775125419245, - 64'd27025025362152, 64'd28493936716347968, - 64'd3814403886660839, 64'd303251651393391, 64'd21028720080409, - 64'd24000428154010, 64'd26566714056631116, - 64'd3888381425628968, 64'd343372202987344, 64'd7413998071180, - 64'd21062492581666, 64'd24611415025440940, - 64'd3927173865649960, 64'd377454151408548, - 64'd5067223338077, - 64'd18225361188348},
		'{64'd4227, 64'd594, - 64'd216, 64'd17, 64'd1, 64'd3992, 64'd561, - 64'd204, 64'd16, 64'd1, 64'd3771, 64'd530, - 64'd192, 64'd15, 64'd1, 64'd3562, 64'd501, - 64'd182, 64'd14, 64'd1, 64'd3364, 64'd473, - 64'd172, 64'd14, 64'd1, 64'd3178, 64'd447, - 64'd162, 64'd13, 64'd1, 64'd3002, 64'd422, - 64'd153, 64'd12, 64'd1, 64'd2835, 64'd399, - 64'd145, 64'd12, 64'd1, 64'd2678, 64'd376, - 64'd137, 64'd11, 64'd1, 64'd2530, 64'd356, - 64'd129, 64'd10, 64'd1, 64'd2390, 64'd336, - 64'd122, 64'd10, 64'd1, 64'd2257, 64'd317, - 64'd115, 64'd9, 64'd1, 64'd2132, 64'd300, - 64'd109, 64'd9, 64'd1, 64'd2014, 64'd283, - 64'd103, 64'd8, 64'd1, 64'd1902, 64'd267, - 64'd97, 64'd8, 64'd0, 64'd1797, 64'd253, - 64'd92, 64'd7, 64'd0, 64'd1697, 64'd239, - 64'd87, 64'd7, 64'd0, 64'd1603, 64'd225, - 64'd82, 64'd7, 64'd0, 64'd1514, 64'd213, - 64'd77, 64'd6, 64'd0, 64'd1430, 64'd201, - 64'd73, 64'd6, 64'd0}};
	localparam logic signed[63:0] Fbr[0:4][0:99] = '{
		'{- 64'd12121701392631576, - 64'd5511085814118572, 64'd179182817565032, 64'd185632095569354, 64'd16375895597195, - 64'd9325598198400832, - 64'd5657779628121171, 64'd40473921396927, 64'd177081116710846, 64'd19110861806506, - 64'd6479371739918228, - 64'd5711846607152701, - 64'd94179714416863, 64'd166074689400989, 64'd21457354306236, - 64'd3628820118258496, - 64'd5675575756494004, - 64'd222828347759746, 64'd152866262543536, 64'd23392124950551, - 64'd818262431874540, - 64'd5552578715388690, - 64'd343681110330425, 64'd137734852169609, 64'd24899090569803, 64'd1910098079483638, - 64'd5347689141144777, - 64'd455128396357463, 64'd120979854632028, 64'd25969340329378, 64'd4516756604170016, - 64'd5066846552975130, - 64'd555760686623897, 64'd102915719072728, 64'd26601031695251, 64'd6965427846254730, - 64'd4716966960170498, - 64'd644383636433401, 64'd83866566471041, 64'd26799180378749, 64'd9223499631869116, - 64'd4305802725520964, - 64'd720029319829657, 64'd64160840461159, 64'd26575351094600, 64'd11262414283044492, - 64'd3841794198979132, - 64'd781963585579850, 64'd44126071739022, 64'd25947257272679, 64'd13057974287534080, - 64'd3333915698514529, - 64'd829689542188433, 64'd24083833356644, 64'd24938278999926, 64'd14590570083431264, - 64'd2791518415715291, - 64'd862947248610265, 64'd4344958634419, 64'd23576909422927, 64'd15845329057963682, - 64'd2224172784336629, - 64'd881709743541835, - 64'd14794913069079, 64'd21896140604860, 64'd16812186111136374, - 64'd1641512772634777, - 64'd886175598422222, - 64'd33059404773208, 64'd19932800397630, 64'd17485877338516620, - 64'd1053084447441928, - 64'd876758226895624, - 64'd50195034455864, 64'd17726852258869, 64'd17865859526355222, - 64'd468201012480347, - 64'd854072225893131, - 64'd65974370219586, 64'd15320670114924, 64'd17956159210960408, 64'd104193651263810, - 64'd818917060201813, - 64'd80198675265970, 64'd12758300349201, 64'd17765156019080896, 64'd655651115491204, - 64'd772258433027506, - 64'd92700018913746, 64'd10084722786950, 64'd17305305865232496, 64'd1178332599016474, - 64'd715207709354171, - 64'd103342838972494, 64'd7345122162380, 64'd16592810325669880, 64'd1665109859989971, - 64'd648999776694870, - 64'd112024949781757, 64'd4584181003857},
		'{- 64'd12121701392629594, - 64'd5511085814118876, 64'd179182817564926, 64'd185632095569345, 64'd16375895597196, - 64'd9325598198398734, - 64'd5657779628121486, 64'd40473921396816, 64'd177081116710836, 64'd19110861806506, - 64'd6479371739916055, - 64'd5711846607153022, - 64'd94179714416977, 64'd166074689400979, 64'd21457354306236, - 64'd3628820118256281, - 64'd5675575756494324, - 64'd222828347759860, 64'd152866262543527, 64'd23392124950551, - 64'd818262431872320, - 64'd5552578715389005, - 64'd343681110330538, 64'd137734852169599, 64'd24899090569804, 64'd1910098079485828, - 64'd5347689141145084, - 64'd455128396357574, 64'd120979854632019, 64'd25969340329379, 64'd4516756604172144, - 64'd5066846552975423, - 64'd555760686624003, 64'd102915719072719, 64'd26601031695252, 64'd6965427846256764, - 64'd4716966960170772, - 64'd644383636433501, 64'd83866566471033, 64'd26799180378749, 64'd9223499631871028, - 64'd4305802725521218, - 64'd720029319829750, 64'd64160840461152, 64'd26575351094601, 64'd11262414283046258, - 64'd3841794198979361, - 64'd781963585579935, 64'd44126071739016, 64'd25947257272679, 64'd13057974287535680, - 64'd3333915698514730, - 64'd829689542188508, 64'd24083833356638, 64'd24938278999926, 64'd14590570083432674, - 64'd2791518415715463, - 64'd862947248610330, 64'd4344958634414, 64'd23576909422928, 64'd15845329057964888, - 64'd2224172784336770, - 64'd881709743541889, - 64'd14794913069083, 64'd21896140604860, 64'd16812186111137364, - 64'd1641512772634885, - 64'd886175598422265, - 64'd33059404773211, 64'd19932800397630, 64'd17485877338517386, - 64'd1053084447442003, - 64'd876758226895655, - 64'd50195034455866, 64'd17726852258869, 64'd17865859526355762, - 64'd468201012480389, - 64'd854072225893150, - 64'd65974370219587, 64'd15320670114924, 64'd17956159210960716, 64'd104193651263801, - 64'd818917060201820, - 64'd80198675265970, 64'd12758300349202, 64'd17765156019080980, 64'd655651115491226, - 64'd772258433027502, - 64'd92700018913746, 64'd10084722786950, 64'd17305305865232360, 64'd1178332599016527, - 64'd715207709354156, - 64'd103342838972492, 64'd7345122162380, 64'd16592810325669532, 64'd1665109859990052, - 64'd648999776694844, - 64'd112024949781754, 64'd4584181003857},
		'{64'd54230251112480224, 64'd10162912064129204, 64'd1107410074232320, 64'd66607254859419, - 64'd34180873857108, 64'd49176792574385560, 64'd10039753153409532, 64'd1154689346203892, 64'd90659314527461, - 64'd27733084614410, 64'd44201062489677208, 64'd9853166970426098, 64'd1189310977363184, 64'd111942322359692, - 64'd21643151376508, 64'd39333038862206016, 64'd9610067924103708, 64'd1212123917937735, 64'd130540713330342, - 64'd15924834974848, 64'd34599287485460208, 64'd9317184474204714, 64'd1223990268590974, 64'd146551387709459, - 64'd10587949604627, 64'd30023063481010368, 64'd8981025649058081, 64'd1225777763232035, 64'd160081907180583, - 64'd5638634772698, 64'd25624428434944856, 64'd8607852106801811, 64'd1218352866297295, 64'd171248769629750, - 64'd1079630659773, 64'd21420380905485056, 64'd8203651557393658, 64'd1202574481872452, 64'd180175768485818, 64'd3089445435503, 64'd17424998170533344, 64'd7774118346376153, 64'd1179288267733101, 64'd186992441354221, 64'd6871823707512, 64'd13649587186875850, 64'd7324636988003550, 64'd1149321543516658, 64'd191832611612620, 64'd10273309452191, 64'd10102842841729462, 64'd6860269424696720, 64'd1113478778790348, 64'd194833025629963, 64'd13302015424023, 64'd6791011690960054, 64'd6385745781726976, 64'd1072537643737978, 64'd196132087331631, 64'd15968100504470, 64'd3718059495358866, 64'd5905458380376236, 64'd1027245602539384, 64'd195868690963791, 64'd18283516061774, 64'd885840985683144, 64'd5423458769409848, 64'd978317027246011, 64'd194181152110122, 64'd20261761204803, - 64'd1705729592333484, 64'd4943457533359528, 64'd926430808047790, 64'd191206236283473, 64'd21917647962927, - 64'd4058508481108936, 64'd4468826636676080, 64'd872228434262854, 64'd187078283753276, 64'd23267077260512, - 64'd6175954170621278, 64'd4002604065104876, 64'd816312519144131, 64'd181928428675371, 64'd24326826399042, - 64'd8062962003819387, 64'd3547500529493366, 64'd759245740666098, 64'd175883910062924, 64'd25114348612645, - 64'd9725702601620356, 64'd3105908002494394, 64'd701550169811212, 64'd169067471673386, 64'd25647585124212, - 64'd11171464967884652, 64'd2679909865120778, 64'd643706957498268, 64'd161596847484811, 64'd25944789999639},
		'{64'd54230251112476992, 64'd10162912064129726, 64'd1107410074232505, 64'd66607254859435, - 64'd34180873857108, 64'd49176792574382072, 64'd10039753153410084, 64'd1154689346204088, 64'd90659314527478, - 64'd27733084614411, 64'd44201062489673520, 64'd9853166970426672, 64'd1189310977363388, 64'd111942322359710, - 64'd21643151376509, 64'd39333038862202176, 64'd9610067924104296, 64'd1212123917937946, 64'd130540713330360, - 64'd15924834974849, 64'd34599287485456248, 64'd9317184474205316, 64'd1223990268591190, 64'd146551387709477, - 64'd10587949604628, 64'd30023063481006344, 64'd8981025649058686, 64'd1225777763232252, 64'd160081907180602, - 64'd5638634772698, 64'd25624428434940792, 64'd8607852106802416, 64'd1218352866297513, 64'd171248769629768, - 64'd1079630659774, 64'd21420380905480984, 64'd8203651557394260, 64'd1202574481872669, 64'd180175768485837, 64'd3089445435502, 64'd17424998170529294, 64'd7774118346376746, 64'd1179288267733315, 64'd186992441354239, 64'd6871823707511, 64'd13649587186871850, 64'd7324636988004131, 64'd1149321543516868, 64'd191832611612637, 64'd10273309452190, 64'd10102842841725546, 64'd6860269424697284, 64'd1113478778790553, 64'd194833025629980, 64'd13302015424022, 64'd6791011690956236, 64'd6385745781727524, 64'd1072537643738176, 64'd196132087331647, 64'd15968100504469, 64'd3718059495355164, 64'd5905458380376764, 64'd1027245602539575, 64'd195868690963806, 64'd18283516061773, 64'd885840985679580, 64'd5423458769410352, 64'd978317027246194, 64'd194181152110136, 64'd20261761204802, - 64'd1705729592336900, 64'd4943457533360008, 64'd926430808047964, 64'd191206236283487, 64'd21917647962926, - 64'd4058508481112190, 64'd4468826636676534, 64'd872228434263020, 64'd187078283753289, 64'd23267077260512, - 64'd6175954170624356, 64'd4002604065105303, 64'd816312519144286, 64'd181928428675384, 64'd24326826399041, - 64'd8062962003822286, 64'd3547500529493765, 64'd759245740666244, 64'd175883910062935, 64'd25114348612645, - 64'd9725702601623068, 64'd3105908002494765, 64'd701550169811348, 64'd169067471673397, 64'd25647585124212, - 64'd11171464967887176, 64'd2679909865121120, 64'd643706957498394, 64'd161596847484821, 64'd25944789999638},
		'{64'd83657983348648656, 64'd9541301882050548, 64'd2521758375897227, 64'd450532855767046, 64'd96732342708448, 64'd79020797936577888, 64'd9012424850491996, 64'd2381976603908496, 64'd425559693579826, 64'd91370441900803, 64'd74640653008692656, 64'd8512863620693828, 64'd2249942974631240, 64'd401970800756419, 64'd86305752754388, 64'd70503300739072888, 64'd8040993209566270, 64'd2125228006348184, 64'd379689446858875, 64'd81521800743706, 64'd66595283062773640, 64'd7595278707286637, 64'd2007426023633749, 64'd358643154638879, 64'd77003024530813, 64'd62903887899153488, 64'd7174270284512957, 64'd1896153837764640, 64'd338763464282259, 64'd72734725347082, 64'd59417107801755872, 64'd6776598476349133, 64'd1791049500275656, 64'd319985710721485, 64'd68703019180740, 64'd56123600900239240, 64'd6400969727721226, 64'd1691771125606240, 64'd302248813291806, 64'd64894791614670, 64'd53012654007306816, 64'd6046162185674793, 64'd1597995779008066, 64'd285495077046799, 64'd61297655167563, 64'd50074147770629656, 64'd5711021724906348, 64'd1509418426096217, 64'd269670005087055, 64'd57899908999662, 64'd47298523756408296, 64'd5394458193600728, 64'd1425750940627034, 64'd254722121291540, 64'd54690500852032, 64'd44676753357501808, 64'd5095441867362750, 64'd1346721167275121, 64'd240602802875004, 64'd51658991095540, 64'd42200308424987944, 64'd4813000099708417, 64'd1272072036360875, 64'd227266122226780, 64'd48795518772615, 64'd39861133527624104, 64'd4546214158220341, 64'd1201560727648924, 64'd214668697516507, 64'd46090769521324, 64'd37651619748974200, 64'd4294216236075956, 64'd1134957880497448, 64'd202769551580809, 64'd43535945277418, 64'd35564579936968036, 64'd4056186629227557, 64'd1072046847789146, 64'd191529978631937, 64'd41122735655812, 64'd33593225325384552, 64'd3831351070052028, 64'd1012622991217009, 64'd180913418354781, 64'd38843290918388, 64'd31731143451212820, 64'd3618978208797132, 64'd956493015632619, 64'd170885336982721, 64'd36690196440209, 64'd29972277296059848, 64'd3418377234631920, 64'd903474340291686, 64'd161413114965480, 64'd34656448591071, 64'd28310905583756036, 64'd3228895628562988, 64'd853394504951638, 64'd152465940863573, 64'd32735431953950}};
	localparam logic signed[63:0] Fbi[0:4][0:99] = '{
		'{- 64'd20467974938558076, 64'd2314420005831342, 64'd1100572195040407, 64'd32611940301810, - 64'd25718338064436, - 64'd21443050477604384, 64'd1584938512519100, 64'd1095333125455362, 64'd54460373751978, - 64'd23086723774012, - 64'd22052921347871056, 64'd855521716972296, 64'd1073297268587196, 64'd74727323968669, - 64'd20186186535086, - 64'd22300465164129556, 64'd137470719399253, 64'd1035373115959941, 64'd93152114409092, - 64'd17070752184426, - 64'd22194077140263000, - 64'd558471004406560, 64'd982684701039992, 64'd109511415021970, - 64'd13795952901513, - 64'd21747353734214364, - 64'd1222265263551204, 64'd916546904696429, 64'd123621442321922, - 64'd10417915813221, - 64'd20978706372071724, - 64'd1844710898556169, 64'd838438636851291, 64'd135339472368277, - 64'd6992473145366, - 64'd19910913597499592, - 64'd2417558109532762, 64'd749974381600231, 64'd144564666397293, - 64'd3574306983146, - 64'd18570620665159952, - 64'd2933604182346382, 64'd652874601994840, 64'd151238219516567, - 64'd216140725251, - 64'd16987796106745588, - 64'd3386769757322648, 64'd548935501598846, 64'd155342853009109, 64'd3032011815140, - 64'd15195155143353004, - 64'd3772155115444260, 64'd439998633116790, 64'd156901680272569, 64'd6123529972295, - 64'd13227559998370616, - 64'd4086076284367489, 64'd327920830212376, 64'd155976485111869, 64'd9015794133221, - 64'd11121407183611766, - 64'd4326081085978768, 64'd214544917552954, 64'd152665458902827, 64'd11670711119996, - 64'd8914011693259571, - 64'd4490945553935468, 64'd101671626696035, 64'd147100449959589, 64'd14055151693393, - 64'd6642997752742528, - 64'd4580651439364955, - 64'd8966887687547, 64'd139443784197307, 64'd16141296364669, - 64'd4345705342420399, - 64'd4596345791716492, - 64'd115731574875758, 64'd129884720830122, 64'd17906887251978, - 64'd2058621160268606, - 64'd4540283846211505, - 64'd217098744416944, 64'd118635610348398, 64'd19335385250248, 64'd183157983446269, - 64'd4415756666453720, - 64'd311679783473965, 64'd105927824362754, 64'd20416033275353, 64'd2346422118907068, - 64'd4227005178100108, - 64'd398238115353751, 64'd92007528088579, 64'd21143827773211, 64'd4400299054528418, - 64'd3979122385158311, - 64'd475703229557823, 64'd77131366294058, 64'd21519402032049},
		'{64'd20467974938559408, - 64'd2314420005831492, - 64'd1100572195040465, - 64'd32611940301814, 64'd25718338064436, 64'd21443050477605440, - 64'd1584938512519208, - 64'd1095333125455406, - 64'd54460373751981, 64'd23086723774012, 64'd22052921347871832, - 64'd855521716972364, - 64'd1073297268587226, - 64'd74727323968671, 64'd20186186535086, 64'd22300465164130044, - 64'd137470719399280, - 64'd1035373115959956, - 64'd93152114409093, 64'd17070752184426, 64'd22194077140263208, 64'd558471004406573, - 64'd982684701039992, - 64'd109511415021970, 64'd13795952901513, 64'd21747353734214296, 64'd1222265263551256, - 64'd916546904696416, - 64'd123621442321920, 64'd10417915813221, 64'd20978706372071392, 64'd1844710898556257, - 64'd838438636851265, - 64'd135339472368274, 64'd6992473145365, 64'd19910913597499008, 64'd2417558109532883, - 64'd749974381600192, - 64'd144564666397289, 64'd3574306983146, 64'd18570620665159136, 64'd2933604182346534, - 64'd652874601994790, - 64'd151238219516562, 64'd216140725251, 64'd16987796106744554, 64'd3386769757322827, - 64'd548935501598786, - 64'd155342853009103, - 64'd3032011815141, 64'd15195155143351782, 64'd3772155115444463, - 64'd439998633116720, - 64'd156901680272563, - 64'd6123529972296, 64'd13227559998369228, 64'd4086076284367710, - 64'd327920830212300, - 64'd155976485111862, - 64'd9015794133222, 64'd11121407183610242, 64'd4326081085979006, - 64'd214544917552871, - 64'd152665458902820, - 64'd11670711119996, 64'd8914011693257937, 64'd4490945553935717, - 64'd101671626695948, - 64'd147100449959581, - 64'd14055151693393, 64'd6642997752740813, 64'd4580651439365210, 64'd8966887687638, - 64'd139443784197299, - 64'd16141296364670, 64'd4345705342418633, 64'd4596345791716750, 64'd115731574875850, - 64'd129884720830115, - 64'd17906887251979, 64'd2058621160266819, 64'd4540283846211762, 64'd217098744417036, - 64'd118635610348390, - 64'd19335385250248, - 64'd183157983448051, 64'd4415756666453972, 64'd311679783474056, - 64'd105927824362747, - 64'd20416033275354, - 64'd2346422118908817, 64'd4227005178100352, 64'd398238115353839, - 64'd92007528088572, - 64'd21143827773212, - 64'd4400299054530106, 64'd3979122385158542, 64'd475703229557907, - 64'd77131366294051, - 64'd21519402032050},
		'{64'd34656575565312940, - 64'd4988108285545681, - 64'd1389538734008945, - 64'd379170625264187, - 64'd67317163494705, 64'd36907080549404824, - 64'd4022832490582728, - 64'd1244312214721891, - 64'd356444177497412, - 64'd66583219400563, 64'd38688484455219192, - 64'd3112083068544692, - 64'd1102567579945230, - 64'd333067760901026, - 64'd65421398079712, 64'd40028568385265104, - 64'd2257829886078850, - 64'd965048182911008, - 64'd309270815359571, - 64'd63877628016734, 64'd40955949332034712, - 64'd1461453472484437, - 64'd832401280626865, - 64'd285265862491704, - 64'd61996651052703, 64'd41499795792327800, - 64'd723786256669338, - 64'd705181638932075, - 64'd261248412089143, - 64'd59821795389116, 64'd41689564127765800, - 64'd45154254508206, - 64'd583855506258482, - 64'd237397002409543, - 64'd57394778848132, 64'd41554755808632264, 64'd574581140706096, - 64'd468804894556953, - 64'd213873362342983, - 64'd54755541201951, 64'd41124695511916016, 64'd1135981582474870, - 64'd360332108951655, - 64'd190822683616961, - 64'd51942104273018, 64'd40428329892898456, 64'd1639990698407458, - 64'd258664470947135, - 64'd168373991424715, - 64'd48990458414845, 64'd39494046712652536, 64'd2087893780182719, - 64'd163959183398814, - 64'd146640602148313, - 64'd45934473909715, 64'd38349513881148224, 64'd2481278467416686, - 64'd76308288930206, - 64'd125720657193185, - 64'd42805835763154, 64'd37021537866946880, 64'd2821996629167747, 64'd4256322993214, - 64'd105697722347071, - 64'd39634000334883, 64'd35535940829298876, 64'd3112127620180786, 64'd77757901573789, - 64'd86641442516250, - 64'd36446172220825, 64'd33917455746356300, 64'd3353943063357565, 64'd144269850470854, - 64'd68608242168432, - 64'd33267299789458, 64'd32189638743641944, 64'd3549873285442806, 64'd203910808051241, - 64'd51642062318009, - 64'd30120087777389, 64'd30374797769297368, 64'd3702475509617544, 64'd256839822823478, - 64'd35775125419248, - 64'd27025025362152, 64'd28493936716348648, 64'd3814403886660708, 64'd303251651393346, - 64'd21028720080413, - 64'd24000428154009, 64'd26566714056631972, 64'd3888381425628816, 64'd343372202987290, - 64'd7413998071185, - 64'd21062492581666, 64'd24611415025441952, 64'd3927173865649788, 64'd377454151408487, 64'd5067223338071, - 64'd18225361188348},
		'{- 64'd34656575565318544, 64'd4988108285546430, 64'd1389538734009220, 64'd379170625264209, 64'd67317163494703, - 64'd36907080549409936, 64'd4022832490583405, 64'd1244312214722141, 64'd356444177497432, 64'd66583219400562, - 64'd38688484455223808, 64'd3112083068545297, 64'd1102567579945454, 64'd333067760901043, 64'd65421398079711, - 64'd40028568385269240, 64'd2257829886079385, 64'd965048182911207, 64'd309270815359586, 64'd63877628016733, - 64'd40955949332038376, 64'd1461453472484904, 64'd832401280627039, 64'd285265862491717, 64'd61996651052702, - 64'd41499795792331008, 64'd723786256669740, 64'd705181638932225, 64'd261248412089155, 64'd59821795389115, - 64'd41689564127768560, 64'd45154254508545, 64'd583855506258609, 64'd237397002409552, 64'd57394778848131, - 64'd41554755808634608, - 64'd574581140705816, 64'd468804894557059, 64'd213873362342991, 64'd54755541201951, - 64'd41124695511917952, - 64'd1135981582474646, 64'd360332108951740, 64'd190822683616967, 64'd51942104273017, - 64'd40428329892900008, - 64'd1639990698407288, 64'd258664470947200, 64'd168373991424719, 64'd48990458414844, - 64'd39494046712653728, - 64'd2087893780182598, 64'd163959183398862, 64'd146640602148316, 64'd45934473909715, - 64'd38349513881149088, - 64'd2481278467416612, 64'd76308288930236, 64'd125720657193187, 64'd42805835763154, - 64'd37021537866947424, - 64'd2821996629167714, - 64'd4256322993199, 64'd105697722347071, 64'd39634000334883, - 64'd35535940829299128, - 64'd3112127620180794, - 64'd77757901573789, 64'd86641442516249, 64'd36446172220825, - 64'd33917455746356280, - 64'd3353943063357609, - 64'd144269850470866, 64'd68608242168430, 64'd33267299789458, - 64'd32189638743641684, - 64'd3549873285442882, - 64'd203910808051266, 64'd51642062318007, 64'd30120087777389, - 64'd30374797769296888, - 64'd3702475509617648, - 64'd256839822823513, 64'd35775125419245, 64'd27025025362152, - 64'd28493936716347968, - 64'd3814403886660839, - 64'd303251651393391, 64'd21028720080409, 64'd24000428154010, - 64'd26566714056631116, - 64'd3888381425628968, - 64'd343372202987344, 64'd7413998071180, 64'd21062492581666, - 64'd24611415025440940, - 64'd3927173865649960, - 64'd377454151408548, - 64'd5067223338077, 64'd18225361188348},
		'{- 64'd4227, 64'd594, 64'd216, 64'd17, - 64'd1, - 64'd3992, 64'd561, 64'd204, 64'd16, - 64'd1, - 64'd3771, 64'd530, 64'd192, 64'd15, - 64'd1, - 64'd3562, 64'd501, 64'd182, 64'd14, - 64'd1, - 64'd3364, 64'd473, 64'd172, 64'd14, - 64'd1, - 64'd3178, 64'd447, 64'd162, 64'd13, - 64'd1, - 64'd3002, 64'd422, 64'd153, 64'd12, - 64'd1, - 64'd2835, 64'd399, 64'd145, 64'd12, - 64'd1, - 64'd2678, 64'd376, 64'd137, 64'd11, - 64'd1, - 64'd2530, 64'd356, 64'd129, 64'd10, - 64'd1, - 64'd2390, 64'd336, 64'd122, 64'd10, - 64'd1, - 64'd2257, 64'd317, 64'd115, 64'd9, - 64'd1, - 64'd2132, 64'd300, 64'd109, 64'd9, - 64'd1, - 64'd2014, 64'd283, 64'd103, 64'd8, - 64'd1, - 64'd1902, 64'd267, 64'd97, 64'd8, - 64'd0, - 64'd1797, 64'd253, 64'd92, 64'd7, - 64'd0, - 64'd1697, 64'd239, 64'd87, 64'd7, - 64'd0, - 64'd1603, 64'd225, 64'd82, 64'd7, - 64'd0, - 64'd1514, 64'd213, 64'd77, 64'd6, - 64'd0, - 64'd1430, 64'd201, 64'd73, 64'd6, - 64'd0}};
	localparam logic signed[63:0] hf[0:1499] = {64'd11691005837312, - 64'd70667902976, - 64'd82071273472, 64'd787514816, 64'd1638997888, 64'd11620470226944, - 64'd211201048576, - 64'd80075431936, 64'd2343618816, 64'd1601011968, 64'd11480201166848, - 64'd349338796032, - 64'd76116705280, 64'd3843500544, 64'd1526184192, 64'd11271788298240, - 64'd483523461120, - 64'd70259892224, 64'd5251344384, 64'd1416697856, 64'd10997584625664, - 64'd612254351360, - 64'd62600273920, 64'd6533577216, 64'd1275646208, 64'd10660677156864, - 64'd734109040640, - 64'd53261762560, 64'd7659540480, 64'd1106893824, 64'd10264840765440, - 64'd847763013632, - 64'd42394480640, 64'd8602073088, 64'd914936320, 64'd9814481567744, - 64'd952008179712, - 64'd30172010496, 64'd9337997312, 64'd704756608, 64'd9314579251200, - 64'd1045768372224, - 64'd16788210688, 64'd9848502272, 64'd481682848, 64'd8770614722560, - 64'd1128113766400, - 64'd2453763840, 64'd10119427072, 64'd251248704, 64'd8188496183296, - 64'd1198272151552, 64'd12607502336, 64'd10141449216, 64'd19058776, 64'd7574474719232, - 64'd1255637778432, 64'd28162451456, 64'd9910159360, - 64'd209339232, 64'd6935062511616, - 64'd1299777847296, 64'd43972554752, 64'd9426054144, - 64'd428573856, 64'd6276944232448, - 64'd1330435850240, 64'd59797811200, 64'd8694424576, - 64'd633559232, 64'd5606887391232, - 64'd1347532488704, 64'd75400634368, 64'd7725167616, - 64'd819593152, 64'd4931656876032, - 64'd1351164100608, 64'd90549592064, 64'd6532513792, - 64'd982442752, 64'd4257923989504, - 64'd1341597810688, 64'd105022963712, 64'd5134683136, - 64'd1118417280, 64'd3592187543552, - 64'd1319265107968, 64'd118612099072, 64'd3553482240, - 64'd1224427008, 64'd2940689973248, - 64'd1284752408576, 64'd131124453376, 64'd1813845120, - 64'd1298028032, 64'd2309344460800, - 64'd1238790045696, 64'd142386298880, - 64'd56666844, - 64'd1337453440, 64'd1703665729536, - 64'd1182239031296, 64'd152245092352, - 64'd2028398464, - 64'd1341629952, 64'd1128708571136, - 64'd1116075982848, 64'd160571424768, - 64'd4070156288, - 64'd1310181248, 64'd589013385216, - 64'd1041377656832, 64'd167260618752, - 64'd6149776384, - 64'd1243418368, 64'd88561303552, - 64'd959302860800, 64'd172233768960, - 64'd8234692608, - 64'd1142317824, - 64'd369263050752, - 64'd871075086336, 64'd175438479360, - 64'd10292500480, - 64'd1008487424, - 64'd781698990080, - 64'd777963503616, 64'd176849125376, - 64'd12291495936, - 64'd844123584, - 64'd1146627948544, - 64'd681264480256, 64'd176466657280, - 64'd14201202688, - 64'd651957504, - 64'd1462582247424, - 64'd582282641408, 64'd174317993984, - 64'd15992844288, - 64'd435194624, - 64'd1728745308160, - 64'd482312617984, 64'd170455089152, - 64'd17639798784, - 64'd197447344, - 64'd1944940969984, - 64'd382621417472, 64'd164953587712, - 64'd19117987840, 64'd57337632, - 64'd2111616581632, - 64'd284431351808, 64'd157911121920, - 64'd20406222848, 64'd324955520, - 64'd2229816000512, - 64'd188904505344, 64'd149445361664, - 64'd21486497792, 64'd601021952, - 64'd2301146169344, - 64'd97128153088, 64'd139691737088, - 64'd22344208384, 64'd881052416, - 64'd2327735959552, - 64'd10101851136, 64'd128801087488, - 64'd22968328192, 64'd1160540928, - 64'd2312190033920, 64'd71273840640, 64'd116936949760, - 64'd23351506944, 64'd1435037312, - 64'd2257536155648, 64'd146206916608, 64'd104272846848, - 64'd23490117632, 64'd1700221056, - 64'd2167170007040, 64'd214021603328, 64'd90989477888, - 64'd23384236032, 64'd1951971072, - 64'd2044793847808, 64'd274164137984, 64'd77271842816, - 64'd23037569024, 64'd2186430208, - 64'd1894356484096, 64'd326206521344, 64'd63306379264, - 64'd22457309184, 64'd2400063744, - 64'd1719988125696, 64'd369848451072, 64'd49278226432, - 64'd21653964800, 64'd2589710848, - 64'd1525937602560, 64'd404917223424, 64'd35368476672, - 64'd20641116160, 64'd2752628480, - 64'd1316508401664, 64'd431365816320, 64'd21751644160, - 64'd19435145216, 64'd2886526976, - 64'd1095996866560, 64'd449269170176, 64'd8593282048, - 64'd18054922240, 64'd2989598208, - 64'd868632363008, 64'd458818879488, - 64'd3952210176, - 64'd16521456640, 64'd3060534528, - 64'd638520852480, 64'd460316344320, - 64'd15743529984, - 64'd14857540608, 64'd3098538240, - 64'd409591775232, 64'd454164316160, - 64'd26654171136, - 64'd13087353856, 64'd3103324416, - 64'd185549750272, 64'd440857657344, - 64'd36573847552, - 64'd11236068352, 64'd3075113728, 64'd30168758272, 64'd420972625920, - 64'd45409632256, - 64'd9329446912, 64'd3014618368, 64'd234433495040, 64'd395155570688, - 64'd53086793728, - 64'd7393442304, 64'd2923020288, 64'd424452390912, 64'd364110905344, - 64'd59549356032, - 64'd5453806592, 64'd2801941504, 64'd597797568512, 64'd328588722176, - 64'd64760328192, - 64'd3535706624, 64'd2653410560, 64'd752424845312, 64'd289372012544, - 64'd68701655040, - 64'd1663370112, 64'd2479820800, 64'd886687268864, 64'd247263887360, - 64'd71373914112, 64'd140252432, 64'd2283885568, 64'd999341621248, 64'd203075092480, - 64'd72795676672, 64'd1853793920, 64'd2068588800, 64'd1089549631488, 64'd157611606016, - 64'd73002688512, 64'd3457744128, 64'd1837133952, 64'd1156872273920, 64'd111662972928, - 64'd72046772224, 64'd4934687232, 64'd1592889088, 64'd1201258758144, 64'd65991131136, - 64'd69994545152, 64'd6269501440, 64'd1339332480, 64'd1223030210560, 64'd21320142848, - 64'd66925940736, 64'd7449516032, 64'd1079996800, 64'd1222858637312, - 64'd21673152512, - 64'd62932586496, 64'd8464630784, 64'd818414592, 64'd1201740447744, - 64'd62367465472, - 64'd58116067328, 64'd9307386880, 64'd558065472, 64'd1160967618560, - 64'd100204232704, - 64'd52586074112, 64'd9973001216, 64'd302324896, 64'd1102094401536, - 64'd134693576704, - 64'd46458503168, 64'd10459357184, 64'd54416568, 64'd1026901737472, - 64'd165419040768, - 64'd39853522944, 64'd10766954496, - 64'd182631840, 64'd937359769600, - 64'd192041009152, - 64'd32893659136, 64'd10898821120, - 64'd406028512, 64'd835588587520, - 64'd214298869760, - 64'd25701863424, 64'd10860393472, - 64'd613252608, 64'd723818905600, - 64'd232011890688, - 64'd18399680512, 64'd10659357696, - 64'd802084352, 64'd604351627264, - 64'd245078786048, - 64'd11105486848, 64'd10305466368, - 64'd970629440, 64'd479518916608, - 64'd253476225024, - 64'd3932826880, 64'd9810327552, - 64'd1117337984, 64'd351645564928, - 64'd257256095744, 64'd3011109376, 64'd9187177472, - 64'd1241017728, 64'd223012421632, - 64'd256541736960, 64'd9626868736, 64'd8450626048, - 64'd1340840704, 64'd95821733888, - 64'd251523268608, 64'd15823948800, 64'd7616397824, - 64'd1416345600, - 64'd27834857472, - 64'd242452021248, 64'd21521836032, 64'd6701065216, - 64'd1467432960, - 64'd146005360640, - 64'd229634211840, 64'd26650853376, 64'd5721768448, - 64'd1494355840, - 64'd256903217152, - 64'd213424111616, 64'd31152828416, 64'd4695947264, - 64'd1497705472, - 64'd358929465344, - 64'd194216591360, 64'd34981539840, 64'd3641068544, - 64'd1478392064, - 64'd450691170304, - 64'd172439420928, 64'd38102986752, 64'd2574366208, - 64'd1437621120, - 64'd531015761920, - 64'd148545306624, 64'd40495456256, 64'd1512592384, - 64'd1376866048, - 64'd598961618944, - 64'd123003813888, 64'd42149396480, 64'd471783904, - 64'd1297838592, - 64'd653824557056, - 64'd96293339136, 64'd43067117568, - 64'd532952512, - 64'd1202454784, - 64'd695139893248, - 64'd68893286400, 64'd43262320640, - 64'd1487633536, - 64'd1092800768, - 64'd722681593856, - 64'd41276420096, 64'd42759462912, - 64'd2379569664, - 64'd971095424, - 64'd736456671232, - 64'd13901696000, 64'd41592975360, - 64'd3197509888, - 64'd839653632, - 64'd736696795136, 64'd12792494080, 64'd39806390272, - 64'd3931759616, - 64'd700848320, - 64'd723846299648, 64'd38394494976, 64'd37451300864, - 64'd4574272000, - 64'd557073088, - 64'd698547699712, 64'd62524903424, 64'd34586300416, - 64'd5118708224, - 64'd410706144, - 64'd661623930880, 64'd84841422848, 64'd31275792384, - 64'd5560475136, - 64'd264074992, - 64'd614059016192, 64'd105042903040, 64'd27588800512, - 64'd5896729088, - 64'd119423504, - 64'd556976635904, 64'd122872651776, 64'd23597715456, - 64'd6126356480, 64'd21118726, - 64'd491616960512, 64'd138120904704, 64'd19377049600, - 64'd6249929728, 64'd155564432, - 64'd419313188864, 64'd150626451456, 64'd15002211328, - 64'd6269634560, 64'd282093536, - 64'd341466644480, 64'd160277495808, 64'd10548287488, - 64'd6189179392, 64'd399074560, - 64'd259522232320, 64'd167011680256, 64'd6088892928, - 64'd6013684224, 64'd505082688, - 64'd174943797248, 64'd170815324160, 64'd1695074048, - 64'd5749549056, 64'd598913920, - 64'd89190154240, 64'd171721965568, - 64'd2565707008, - 64'd5404309504, 64'd679595200, - 64'd3691991296, 64'd169810132992, - 64'd6630496768, - 64'd4986481152, 64'd746391296, 64'd80169967616, 64'd165200642048, - 64'd10441671680, - 64'd4505391104, 64'd798807168, 64'd161085259776, 64'd158053154816, - 64'd13947649024, - 64'd3971005440, 64'd836586944, 64'd237832192000, 64'd148562329600, - 64'd17103477760, - 64'd3393752832, 64'd859709248, 64'd309294268416, 64'd136953618432, - 64'd19871305728, - 64'd2784346368, 64'd868379008, 64'd374474440704, 64'd123478548480, - 64'd22220722176, - 64'd2153606912, 64'd863016384, 64'd432506929152, 64'd108409978880, - 64'd24128972800, - 64'd1512292864, 64'd844242304, 64'd482666741760, 64'd92037005312, - 64'd25581041664, - 64'd870935104, 64'd812862080, 64'd524376375296, 64'd74659897344, - 64'd26569621504, - 64'd239681664, 64'd769845952, 64'd557210140672, 64'd56584978432, - 64'd27094951936, 64'd371845536, 64'd716308672, 64'd580896161792, 64'd38119600128, - 64'd27164561408, 64'd954681536, 64'd653486912, 64'd595315195904, 64'd19567282176, - 64'd26792882176, 64'd1500634240, 64'd582715968, 64'd600498044928, 64'd1223063168, - 64'd26000803840, 64'd2002384256, 64'd505405504, 64'd596619952128, - 64'd16630842368, - 64'd24815104000, 64'd2453567488, 64'd423015232, 64'd583993196544, - 64'd33729054720, - 64'd23267842048, 64'd2848840704, 64'd337030624, 64'd563057786880, - 64'd49826627584, - 64'd21395662848, 64'd3183928064, 64'd248938832, 64'd534370353152, - 64'd64702210048, - 64'd19239073792, 64'd3455651072, 64'd160205840, 64'd498591858688, - 64'd78160740352, - 64'd16841673728, 64'd3661937664, 64'd72254360, 64'd456473706496, - 64'd90035634176, - 64'd14249368576, 64'd3801817344, - 64'd13556562, 64'd408843091968, - 64'd100190420992, - 64'd11509573632, 64'd3875396352, - 64'd95950400, 64'd356587700224, - 64'd108519923712, - 64'd8670417920, 64'd3883819008, - 64'd173750016, 64'd300639846400, - 64'd114950856704, - 64'd5779971072, 64'd3829213440, - 64'd245892384, 64'd241960419328, - 64'd119441907712, - 64'd2885491200, 64'd3714623232, - 64'd311441088, 64'd181523120128, - 64'd121983336448, - 64'd32715716, 64'd3543929344, - 64'd369596384, 64'd120298782720, - 64'd122596114432, 64'd2734803712, 64'd3321759488, - 64'd419702784, 64'd59240333312, - 64'd121330532352, 64'd5376306176, 64'd3053389312, - 64'd461254144, - 64'd731416192, - 64'd118264520704, 64'd7854364160, 64'd2744639488, - 64'd493896352, - 64'd58741088256, - 64'd113501454336, 64'd10135356416, 64'd2401764352, - 64'd517427488, - 64'd113970864128, - 64'd107167793152, 64'd12189862912, 64'd2031339264, - 64'd531795584, - 64'd165671337984, - 64'd99410255872, 64'd13992983552, 64'd1640147840, - 64'd537094144, - 64'd213170946048, - 64'd90392961024, 64'd15524575232, 64'd1235068032, - 64'd533555648, - 64'd255883870208, - 64'd80294240256, 64'd16769404928, 64'd822961600, - 64'd521543200, - 64'd293316329472, - 64'd69303451648, 64'd17717221376, 64'd410567744, - 64'd501540064, - 64'd325071339520, - 64'd57617629184, 64'd18362755072, 64'd4401630, - 64'd474138144, - 64'd350851596288, - 64'd45438197760, 64'd18705618944, - 64'd389339424, - 64'd440024864, - 64'd370460917760, - 64'd32967698432, 64'd18750169088, - 64'd764861952, - 64'd399969216, - 64'd383804112896, - 64'd20406595584, 64'd18505261056, - 64'd1116853120, - 64'd354806880, - 64'd390884950016, - 64'd7950255616, 64'd17983975424, - 64'd1440547328, - 64'd305424896, - 64'd391803043840, 64'd4213928448, 64'd17203263488, - 64'd1731781888, - 64'd252746048, - 64'd386749202432, 64'd15909174272, 64'd16183558144, - 64'd1987041664, - 64'd197713280, - 64'd375999365120, 64'd26971701248, 64'd14948338688, - 64'd2203492096, - 64'd141274192, - 64'd359907786752, 64'd37252841472, 64'd13523662848, - 64'd2379000320, - 64'd84366160, - 64'd338898780160, 64'd46620835840, 64'd11937680384, - 64'd2512144384, - 64'd27902050, - 64'd313458130944, 64'd54962319360, 64'd10220119040, - 64'd2602212096, 64'd27243218, - 64'd284123299840, 64'd62183481344, 64'd8401773568, - 64'd2649188096, 64'd80245000, - 64'd251473739776, 64'd68210851840, 64'd6513990144, - 64'd2653730304, 64'd130340104, - 64'd216120344576, 64'd72991768576, 64'd4588161536, - 64'd2617136384, 64'd176836592, - 64'd178695159808, 64'd76494503936, 64'd2655238656, - 64'd2541304064, 64'd219122144, - 64'd139840864256, 64'd78708088832, 64'd745262912, - 64'd2428679424, 64'd256670928, - 64'd100200562688, 64'd79641739264, - 64'd1113069184, - 64'd2282201088, 64'd289048864, - 64'd60407840768, 64'd79324094464, - 64'd2892806656, - 64'd2105238400, 64'd315917216, - 64'd21077354496, 64'd77802110976, - 64'd4569103872, - 64'd1901523584, 64'd337034816, 64'd17204037632, 64'd75139710976, - 64'd6119537152, - 64'd1675082368, 64'd352258336, 64'd53885362176, 64'd71416266752, - 64'd7524370432, - 64'd1430161280, 64'd361541280, 64'd88458821632, 64'd66724818944, - 64'd8766772224, - 64'd1171153920, 64'd364931584, 64'd120466178048, 64'd61170216960, - 64'd9832982528, - 64'd902527872, 64'd362567392, 64'd149504163840, 64'd54867099648, - 64'd10712419328, - 64'd628753024, 64'd354672160, 64'd175228796928, 64'd47937769472, - 64'd11397739520, - 64'd354231488, 64'd341548192, 64'd197358780416, 64'd40510091264, - 64'd11884845056, - 64'd83231856, 64'd323569152, 64'd215677616128, 64'd32715292672, - 64'd12172835840, 64'd180172848, 64'd301172096, 64'd230034898944, 64'd24685850624, - 64'd12263920640, 64'd432161888, 64'd274848320, 64'd240346251264, 64'd16553392128, - 64'd12163275776, 64'd669217728, 64'd245134048, 64'd246592552960, 64'd8446690816, - 64'd11878867968, 64'd888170560, 64'd212600496, 64'd248817893376, 64'd489775968, - 64'd11421236224, 64'd1086235904, 64'd177843856, 64'd247126884352, - 64'd7199825408, - 64'd10803245056, 64'd1261044992, 64'd141475104, 64'd241680891904, - 64'd14512684032, - 64'd10039804928, 64'd1410667520, 64'd104110152, 64'd232693678080, - 64'd21348886528, - 64'd9147576320, 64'd1533627520, 64'd66359960, 64'd220426354688, - 64'd27619258368, - 64'd8144650752, 64'd1628909952, 64'd28821298, 64'd205181698048, - 64'd33246382080, - 64'd7050222080, 64'd1695962624, - 64'd7932100, 64'd187298070528, - 64'd38165393408, - 64'd5884255744, 64'd1734687744, - 64'd43357656, 64'd167143030784, - 64'd42324561920, - 64'd4667152384, 64'd1745429632, - 64'd76951352, 64'd145106616320, - 64'd45685649408, - 64'd3419417088, 64'd1728953472, - 64'd108254256, 64'd121594593280, - 64'd48224038912, - 64'd2161339904, 64'd1686420352, - 64'd136858144, 64'd97021640704, - 64'd49928663040, - 64'd912688192, 64'd1619355392, - 64'd162410176, 64'd71804624896, - 64'd50801717248, 64'd307581728, 64'd1529612416, - 64'd184616448, 64'd46356127744, - 64'd50858168320, 64'd1481589760, 64'd1419333760, - 64'd203244672, 64'd21078155264, - 64'd50125090816, 64'd2592772864, 64'd1290908032, - 64'd218125648, - 64'd3643667456, - 64'd48640860160, 64'd3626097664, 64'd1146924288, - 64'd229153872, - 64'd27445524480, - 64'd46454153216, 64'd4568240128, 64'd990125760, - 64'd236286912, - 64'd49990291456, - 64'd43622846464, 64'd5407735808, 64'd823361984, - 64'd239544096, - 64'd70971834368, - 64'd40212836352, 64'd6135093248, 64'd649540928, - 64'd239004064, - 64'd90118692864, - 64'd36296716288, 64'd6742875648, 64'd471582400, - 64'd234801584, - 64'd107197112320, - 64'd31952439296, 64'd7225745408, 64'd292372320, - 64'd227123632, - 64'd122013368320, - 64'd27261941760, 64'd7580477440, 64'd114718976, - 64'd216204656, - 64'd134415384576, - 64'd22309724160, 64'd7805936128, - 64'd58687512, - 64'd202321472, - 64'd144293707776, - 64'd17181462528, 64'd7903024128, - 64'd225313088, - 64'd185787472, - 64'd151581720576, - 64'd11962642432, 64'd7874598400, - 64'd382813664, - 64'd166946560, - 64'd156255223808, - 64'd6737245696, 64'd7725361664, - 64'd529064992, - 64'd146166848, - 64'd158331387904, - 64'd1586496384, 64'd7461724672, - 64'd662188224, - 64'd123834096, - 64'd157867048960, 64'd3412300288, 64'd7091653120, - 64'd780570624, - 64'd100345176, - 64'd154956480512, 64'd8186822656, 64'd6624487424, - 64'd882881728, - 64'd76101528, - 64'd149728690176, 64'd12670684160, 64'd6070755840, - 64'd968084352, - 64'd51502828, - 64'd142344208384, 64'd16804258816, 64'd5441968640, - 64'd1035440832, - 64'd26940826, - 64'd132991549440, 64'd20535373824, 64'd4750409216, - 64'd1084514176, - 64'd2793569, - 64'd121883320320, 64'd23819872256, 64'd4008914176, - 64'd1115165056, 64'd20580006, - 64'd109252124672, 64'd26622011392, 64'd3230659840, - 64'd1127543552, 64'd42844976, - 64'd95346270208, 64'd28914745344, 64'd2428945152, - 64'd1122077440, 64'd63694820, - 64'd80425385984, 64'd30679842816, 64'd1616980608, - 64'd1099455744, 64'd82855200, - 64'd64756006912, 64'd31907868672, 64'd807688704, - 64'd1060610112, 64'd100087128, - 64'd48607227904, 64'd32598034432, 64'd13512165, - 64'd1006691072, 64'd115189488, - 64'd32246421504, 64'd32757919744, - 64'd753761856, - 64'd939043776, 64'd128000856, - 64'd15935166464, 64'd32403066880, - 64'd1483162240, - 64'd859180288, 64'd138400672, 64'd74618512, 64'd31556468736, - 64'd2164676096, - 64'd768750464, 64'd146309760, 64'd15544250368, 64'd30247966720, - 64'd2789371904, - 64'd669511808, 64'd151690080, 64'd30251536384, 64'd28513552384, - 64'd3349500416, - 64'd563298944, 64'd154544048, 64'd43993653248, 64'd26394601472, - 64'd3838575360, - 64'd451992000, 64'd154913040, 64'd56589647872, 64'd23937046528, - 64'd4251430912, - 64'd337486560, 64'd152875456, 64'd67882487808, 64'd21190518784, - 64'd4584256512, - 64'd221663488, 64'd148544336, 64'd77740703744, 64'd18207447040, - 64'd4834612224, - 64'd106360376, 64'd142064320, 64'd86059532288, 64'd15042149376, - 64'd5001415680, 64'd6655432, 64'd133608432, 64'd92761669632, 64'd11749935104, - 64'd5084918784, 64'd115711832, 64'd123374440, 64'd97797521408, 64'd8386205184, - 64'd5086653952, 64'd219254640, 64'd111580928, 64'd101145042944, 64'd5005594624, - 64'd5009368576, 64'd315867680, 64'd98463200, 64'd102809133056, 64'd1661150336, - 64'd4856942592, 64'd404289984, 64'd84269136, 64'd102820667392, - 64'd1596436608, - 64'd4634288128, 64'd483430176, 64'd69254864, 64'd101235122176, - 64'd4719538176, - 64'd4347238912, 64'd552377600, 64'd53680552, 64'd98130878464, - 64'd7664223744, - 64'd4002430464, 64'd610410112, 64'd37806244, 64'd93607264256, - 64'd10390815744, - 64'd3607167488, 64'd656999424, 64'd21887816, 64'd87782260736, - 64'd12864362496, - 64'd3169290496, 64'd691811968, 64'd6173181, 64'd80790077440, - 64'd15055016960, - 64'd2697033984, 64'd714708224, - 64'd9101296, 64'd72778498048, - 64'd16938331136, - 64'd2198887424, 64'd725737856, - 64'd23714064, 64'd63906152448, - 64'd18495447040, - 64'd1683453824, 64'd725132608, - 64'd37461312, 64'd54339653632, - 64'd19713210368, - 64'd1159312768, 64'd713296768, - 64'd50159536, 64'd44250787840, - 64'd20584165376, - 64'd634889024, 64'd690794752, - 64'd61647676, 64'd33813639168, - 64'd21106491392, - 64'd118326248, 64'd658337280, - 64'd71788872, 64'd23201835008, - 64'd21283842048, 64'd382629120, 64'd616765184, - 64'd80471752, 64'd12585860096, - 64'd21125087232, 64'd860734720, 64'd567032064, - 64'd87611304, 64'd2130512896, - 64'd20644018176, 64'd1309347456, 64'd510185696, - 64'd93149288, - 64'd8007448576, - 64'd19858956288, 64'd1722505984, 64'd447348576, - 64'd97054256, - 64'd17681471488, - 64'd18792316928, 64'd2095000448, 64'd379698048, - 64'd99321104, - 64'd26757134336, - 64'd17470130176, 64'd2422427648, 64'd308446240, - 64'd99970280, - 64'd35113828352, - 64'd15921509376, 64'd2701231360, 64'd234820016, - 64'd99046608, - 64'd42646147072, - 64'd14178094080, 64'd2928730368, 64'd160041504, - 64'd96617760, - 64'd49265025024, - 64'd12273478656, 64'd3103128832, 64'd85309368, - 64'd92772416, - 64'd54898561024, - 64'd10242625536, 64'd3223515136, 64'd11780941, - 64'd87618232, - 64'd59492548608, - 64'd8121272832, 64'd3289845760, - 64'd59444232, - 64'd81279464, - 64'd63010721792, - 64'd5945358336, 64'd3302916864, - 64'd127339528, - 64'd73894544, - 64'd65434730496, - 64'd3750452736, 64'd3264323072, - 64'd190964656, - 64'd65613412, - 64'd66763780096, - 64'd1571222144, 64'd3176407040, - 64'd249477360, - 64'd56594828, - 64'd67014103040, 64'd559078976, 64'd3042195712, - 64'd302143104, - 64'd47003604, - 64'd66218090496, 64'd2609076224, 64'd2865332736, - 64'd348342816, - 64'd37007848, - 64'd64423264256, 64'd4549698048, 64'd2649999360, - 64'd387578592, - 64'd26776244, - 64'd61691031552, 64'd6354548224, 64'd2400832000, - 64'd419477408, - 64'd16475429, - 64'd58095259648, 64'd8000225280, 64'd2122835328, - 64'd443792480, - 64'd6267468, - 64'd53720711168, 64'd9466584064, 64'd1821291904, - 64'd460403008, 64'd3692493, - 64'd48661364736, 64'd10736937984, 64'd1501670912, - 64'd469311648, 64'd13258402, - 64'd43018645504, 64'd11798201344, 64'd1169537280, - 64'd470640448, 64'd22295256, - 64'd36899602432, 64'd12640969728, 64'd830462080, - 64'd464624800, 64'd30680818, - 64'd30415069184, 64'd13259542528, 64'd489935872, - 64'd451606016, 64'd38307084, - 64'd23677794304, 64'd13651887104, 64'd153286496, - 64'd432022368, 64'd45081468, - 64'd16800658432, 64'd13819544576, - 64'd174398144, - 64'd406399232, 64'd50927724, - 64'd9894899712, 64'd13767486464, - 64'd488340800, - 64'd375337760, 64'd55786572, - 64'd3068452864, 64'd13503922176, - 64'd784138432, - 64'd339503104, 64'd59616036, 64'd3575611392, 64'd13040061440, - 64'd1057817792, - 64'd299612032, 64'd62391524, 64'd9940521984, 64'd12389841920, - 64'd1305882624, - 64'd256419936, 64'd64105612, 64'd15937092608, 64'd11569616896, - 64'd1525351552, - 64'd210707840, 64'd64767576, 64'd21484853248, 64'd10597824512, - 64'd1713787136, - 64'd163269520, 64'd64402692, 64'd26512994304, 64'd9494629376, - 64'd1869315200, - 64'd114898680, 64'd63051300, 64'd30961149952, 64'd8281552384, - 64'd1990634752, - 64'd66376692, 64'd60767672, 64'd34779967488, 64'd6981092352, - 64'd2077019008, - 64'd18460890, 64'd57618692, 64'd37931511808, 64'd5616342528, - 64'd2128306816, 64'd28126356, 64'd53682408, 64'd40389468160, 64'd4210614016, - 64'd2144887040, 64'd72707656, 64'd49046428, 64'd42139148288, 64'd2787066880, - 64'd2127672832, 64'd114659568, 64'd43806252, 64'd43177336832, 64'd1368355968, - 64'd2078070528, 64'd153420464, 64'd38063520, 64'd43511943168, - 64'd23702650, - 64'd1997940864, 64'd188497136, 64'd31924228, 64'd43161522176, - 64'd1368441600, - 64'd1889554944, 64'd219470112, 64'd25496940, 64'd42154598400, - 64'd2646623744, - 64'd1755545344, 64'd245997696, 64'd18891022, 64'd40528924672, - 64'd3840692224, - 64'd1598852736, 64'd267818624, 64'd12214913, 64'd38330544128, - 64'd4934985728, - 64'd1422670208, 64'd284753408, 64'd5574480, 64'd35612844032, - 64'd5915916800, - 64'd1230385152, 64'd296704352, - 64'd928537, 64'd32435431424, - 64'd6772112896, - 64'd1025520192, 64'd303654304, - 64'd7197964, 64'd28863043584, - 64'd7494518784, - 64'd811674048, 64'd305664192, - 64'd13144493, 64'd24964341760, - 64'd8076455424, - 64'd592463360, 64'd302869440, - 64'd18686836, 64'd20810729472, - 64'd8513648640, - 64'd371465760, 64'd295475424, - 64'd23752716, 64'd16475149312, - 64'd8804207616, - 64'd152165872, 64'd283751840, - 64'd28279676, 64'd12030904320, - 64'd8948580352, 64'd62095476, 64'd268026352, - 64'd32215728, 64'd7550502912, - 64'd8949464064, 64'd268168304, 64'd248677680, - 64'd35519788, 64'd3104569856, - 64'd8811685888, 64'd463135744, 64'd226127840, - 64'd38161968, - 64'd1239189120, - 64'd8542060544, 64'd644351488, 64'd200834240, - 64'd40123628, - 64'd5416935936, - 64'd8149216256, 64'd809471616, 64'd173281424, - 64'd41397324, - 64'd9369559040, - 64'd7643397120, 64'd956480640, 64'd143972544, - 64'd41986520, - 64'd13043429376, - 64'd7036254208, 64'd1083711744, 64'd113421008, - 64'd41905164, - 64'd16391049216, - 64'd6340613120, 64'd1189860736, 64'd82142176, - 64'd41177136, - 64'd19371575296, - 64'd5570238976, 64'd1273994496, 64'd50645276, - 64'd39835528, - 64'd21951229952, - 64'd4739590656, 64'd1335551872, 64'd19425748, - 64'd37921832, - 64'd24103593984, - 64'd3863571968, 64'd1374341120, - 64'd11041996, - 64'd35484996, - 64'd25809750016, - 64'd2957286656, 64'd1390529536, - 64'd40311192, - 64'd32580432, - 64'd27058341888, - 64'd2035798272, 64'd1384628608, - 64'd67968728, - 64'd29268928, - 64'd27845476352, - 64'd1113897088, 64'd1357475456, - 64'd93640400, - 64'd25615532, - 64'd28174551040, - 64'd205880560, 64'd1310208000, - 64'd116995408, - 64'd21688388, - 64'd28055937024, 64'd674651648, 64'd1244237184, - 64'd137750016, - 64'd17557590, - 64'd27506599936, 64'd1514984704, 64'd1161216512, - 64'd155670336, - 64'd13294021, - 64'd26549600256, 64'd2303456000, 64'd1063007808, - 64'd170574336, - 64'd8968230, - 64'd25213538304, 64'd3029600256, 64'd951645312, - 64'd182332832, - 64'd4649348, - 64'd23531919360, 64'd3684270848, 64'd829298368, - 64'd190869744, - 64'd404071, - 64'd21542475776, 64'd4259737856, 64'd698233472, - 64'd196161488, 64'd3704301, - 64'd19286431744, 64'd4749759488, 64'd560775680, - 64'd198235584, 64'd7616722, - 64'd16807752704, 64'd5149628416, 64'd419270496, - 64'd197168432, 64'd11279177, - 64'd14152366080, 64'd5456193024, 64'd276047136, - 64'd193082576, 64'd14643346, - 64'd11367388160, 64'd5667854336, 64'd133382744, - 64'd186143184, 64'd17667162, - 64'd8500353536, 64'd5784537600, - 64'd6531030, - 64'd176554064, 64'd20315252, - 64'd5598459904, 64'd5807642112, - 64'd141619152, - 64'd164553216, 64'd22559258, - 64'd2707853312, 64'd5739970048, - 64'd269951392, - 64'd150407984, 64'd24378042, 64'd127054280, 64'd5585635840, - 64'd389767392, - 64'd134409888, 64'd25757768, 64'd2864213504, 64'd5349958144, - 64'd499498080, - 64'd116869344, 64'd26691872, 64'd5464509952, 64'd5039334912, - 64'd597783744, - 64'd98110200, 64'd27180914};
	localparam logic signed[63:0] hb[0:1499] = {64'd11691005837312, 64'd70667902976, - 64'd82071273472, - 64'd787514816, 64'd1638997888, 64'd11620470226944, 64'd211201048576, - 64'd80075431936, - 64'd2343618816, 64'd1601011968, 64'd11480201166848, 64'd349338796032, - 64'd76116705280, - 64'd3843500544, 64'd1526184192, 64'd11271788298240, 64'd483523461120, - 64'd70259892224, - 64'd5251344384, 64'd1416697856, 64'd10997584625664, 64'd612254351360, - 64'd62600273920, - 64'd6533577216, 64'd1275646208, 64'd10660677156864, 64'd734109040640, - 64'd53261762560, - 64'd7659540480, 64'd1106893824, 64'd10264840765440, 64'd847763013632, - 64'd42394480640, - 64'd8602073088, 64'd914936320, 64'd9814481567744, 64'd952008179712, - 64'd30172010496, - 64'd9337997312, 64'd704756608, 64'd9314579251200, 64'd1045768372224, - 64'd16788210688, - 64'd9848502272, 64'd481682848, 64'd8770614722560, 64'd1128113766400, - 64'd2453763840, - 64'd10119427072, 64'd251248704, 64'd8188496183296, 64'd1198272151552, 64'd12607502336, - 64'd10141449216, 64'd19058776, 64'd7574474719232, 64'd1255637778432, 64'd28162451456, - 64'd9910159360, - 64'd209339232, 64'd6935062511616, 64'd1299777847296, 64'd43972554752, - 64'd9426054144, - 64'd428573856, 64'd6276944232448, 64'd1330435850240, 64'd59797811200, - 64'd8694424576, - 64'd633559232, 64'd5606887391232, 64'd1347532488704, 64'd75400634368, - 64'd7725167616, - 64'd819593152, 64'd4931656876032, 64'd1351164100608, 64'd90549592064, - 64'd6532513792, - 64'd982442752, 64'd4257923989504, 64'd1341597810688, 64'd105022963712, - 64'd5134683136, - 64'd1118417280, 64'd3592187543552, 64'd1319265107968, 64'd118612099072, - 64'd3553482240, - 64'd1224427008, 64'd2940689973248, 64'd1284752408576, 64'd131124453376, - 64'd1813845120, - 64'd1298028032, 64'd2309344460800, 64'd1238790045696, 64'd142386298880, 64'd56666844, - 64'd1337453440, 64'd1703665729536, 64'd1182239031296, 64'd152245092352, 64'd2028398464, - 64'd1341629952, 64'd1128708571136, 64'd1116075982848, 64'd160571424768, 64'd4070156288, - 64'd1310181248, 64'd589013385216, 64'd1041377656832, 64'd167260618752, 64'd6149776384, - 64'd1243418368, 64'd88561303552, 64'd959302860800, 64'd172233768960, 64'd8234692608, - 64'd1142317824, - 64'd369263050752, 64'd871075086336, 64'd175438479360, 64'd10292500480, - 64'd1008487424, - 64'd781698990080, 64'd777963503616, 64'd176849125376, 64'd12291495936, - 64'd844123584, - 64'd1146627948544, 64'd681264480256, 64'd176466657280, 64'd14201202688, - 64'd651957504, - 64'd1462582247424, 64'd582282641408, 64'd174317993984, 64'd15992844288, - 64'd435194624, - 64'd1728745308160, 64'd482312617984, 64'd170455089152, 64'd17639798784, - 64'd197447344, - 64'd1944940969984, 64'd382621417472, 64'd164953587712, 64'd19117987840, 64'd57337632, - 64'd2111616581632, 64'd284431351808, 64'd157911121920, 64'd20406222848, 64'd324955520, - 64'd2229816000512, 64'd188904505344, 64'd149445361664, 64'd21486497792, 64'd601021952, - 64'd2301146169344, 64'd97128153088, 64'd139691737088, 64'd22344208384, 64'd881052416, - 64'd2327735959552, 64'd10101851136, 64'd128801087488, 64'd22968328192, 64'd1160540928, - 64'd2312190033920, - 64'd71273840640, 64'd116936949760, 64'd23351506944, 64'd1435037312, - 64'd2257536155648, - 64'd146206916608, 64'd104272846848, 64'd23490117632, 64'd1700221056, - 64'd2167170007040, - 64'd214021603328, 64'd90989477888, 64'd23384236032, 64'd1951971072, - 64'd2044793847808, - 64'd274164137984, 64'd77271842816, 64'd23037569024, 64'd2186430208, - 64'd1894356484096, - 64'd326206521344, 64'd63306379264, 64'd22457309184, 64'd2400063744, - 64'd1719988125696, - 64'd369848451072, 64'd49278226432, 64'd21653964800, 64'd2589710848, - 64'd1525937602560, - 64'd404917223424, 64'd35368476672, 64'd20641116160, 64'd2752628480, - 64'd1316508401664, - 64'd431365816320, 64'd21751644160, 64'd19435145216, 64'd2886526976, - 64'd1095996866560, - 64'd449269170176, 64'd8593282048, 64'd18054922240, 64'd2989598208, - 64'd868632363008, - 64'd458818879488, - 64'd3952210176, 64'd16521456640, 64'd3060534528, - 64'd638520852480, - 64'd460316344320, - 64'd15743529984, 64'd14857540608, 64'd3098538240, - 64'd409591775232, - 64'd454164316160, - 64'd26654171136, 64'd13087353856, 64'd3103324416, - 64'd185549750272, - 64'd440857657344, - 64'd36573847552, 64'd11236068352, 64'd3075113728, 64'd30168758272, - 64'd420972625920, - 64'd45409632256, 64'd9329446912, 64'd3014618368, 64'd234433495040, - 64'd395155570688, - 64'd53086793728, 64'd7393442304, 64'd2923020288, 64'd424452390912, - 64'd364110905344, - 64'd59549356032, 64'd5453806592, 64'd2801941504, 64'd597797568512, - 64'd328588722176, - 64'd64760328192, 64'd3535706624, 64'd2653410560, 64'd752424845312, - 64'd289372012544, - 64'd68701655040, 64'd1663370112, 64'd2479820800, 64'd886687268864, - 64'd247263887360, - 64'd71373914112, - 64'd140252432, 64'd2283885568, 64'd999341621248, - 64'd203075092480, - 64'd72795676672, - 64'd1853793920, 64'd2068588800, 64'd1089549631488, - 64'd157611606016, - 64'd73002688512, - 64'd3457744128, 64'd1837133952, 64'd1156872273920, - 64'd111662972928, - 64'd72046772224, - 64'd4934687232, 64'd1592889088, 64'd1201258758144, - 64'd65991131136, - 64'd69994545152, - 64'd6269501440, 64'd1339332480, 64'd1223030210560, - 64'd21320142848, - 64'd66925940736, - 64'd7449516032, 64'd1079996800, 64'd1222858637312, 64'd21673152512, - 64'd62932586496, - 64'd8464630784, 64'd818414592, 64'd1201740447744, 64'd62367465472, - 64'd58116067328, - 64'd9307386880, 64'd558065472, 64'd1160967618560, 64'd100204232704, - 64'd52586074112, - 64'd9973001216, 64'd302324896, 64'd1102094401536, 64'd134693576704, - 64'd46458503168, - 64'd10459357184, 64'd54416568, 64'd1026901737472, 64'd165419040768, - 64'd39853522944, - 64'd10766954496, - 64'd182631840, 64'd937359769600, 64'd192041009152, - 64'd32893659136, - 64'd10898821120, - 64'd406028512, 64'd835588587520, 64'd214298869760, - 64'd25701863424, - 64'd10860393472, - 64'd613252608, 64'd723818905600, 64'd232011890688, - 64'd18399680512, - 64'd10659357696, - 64'd802084352, 64'd604351627264, 64'd245078786048, - 64'd11105486848, - 64'd10305466368, - 64'd970629440, 64'd479518916608, 64'd253476225024, - 64'd3932826880, - 64'd9810327552, - 64'd1117337984, 64'd351645564928, 64'd257256095744, 64'd3011109376, - 64'd9187177472, - 64'd1241017728, 64'd223012421632, 64'd256541736960, 64'd9626868736, - 64'd8450626048, - 64'd1340840704, 64'd95821733888, 64'd251523268608, 64'd15823948800, - 64'd7616397824, - 64'd1416345600, - 64'd27834857472, 64'd242452021248, 64'd21521836032, - 64'd6701065216, - 64'd1467432960, - 64'd146005360640, 64'd229634211840, 64'd26650853376, - 64'd5721768448, - 64'd1494355840, - 64'd256903217152, 64'd213424111616, 64'd31152828416, - 64'd4695947264, - 64'd1497705472, - 64'd358929465344, 64'd194216591360, 64'd34981539840, - 64'd3641068544, - 64'd1478392064, - 64'd450691170304, 64'd172439420928, 64'd38102986752, - 64'd2574366208, - 64'd1437621120, - 64'd531015761920, 64'd148545306624, 64'd40495456256, - 64'd1512592384, - 64'd1376866048, - 64'd598961618944, 64'd123003813888, 64'd42149396480, - 64'd471783904, - 64'd1297838592, - 64'd653824557056, 64'd96293339136, 64'd43067117568, 64'd532952512, - 64'd1202454784, - 64'd695139893248, 64'd68893286400, 64'd43262320640, 64'd1487633536, - 64'd1092800768, - 64'd722681593856, 64'd41276420096, 64'd42759462912, 64'd2379569664, - 64'd971095424, - 64'd736456671232, 64'd13901696000, 64'd41592975360, 64'd3197509888, - 64'd839653632, - 64'd736696795136, - 64'd12792494080, 64'd39806390272, 64'd3931759616, - 64'd700848320, - 64'd723846299648, - 64'd38394494976, 64'd37451300864, 64'd4574272000, - 64'd557073088, - 64'd698547699712, - 64'd62524903424, 64'd34586300416, 64'd5118708224, - 64'd410706144, - 64'd661623930880, - 64'd84841422848, 64'd31275792384, 64'd5560475136, - 64'd264074992, - 64'd614059016192, - 64'd105042903040, 64'd27588800512, 64'd5896729088, - 64'd119423504, - 64'd556976635904, - 64'd122872651776, 64'd23597715456, 64'd6126356480, 64'd21118726, - 64'd491616960512, - 64'd138120904704, 64'd19377049600, 64'd6249929728, 64'd155564432, - 64'd419313188864, - 64'd150626451456, 64'd15002211328, 64'd6269634560, 64'd282093536, - 64'd341466644480, - 64'd160277495808, 64'd10548287488, 64'd6189179392, 64'd399074560, - 64'd259522232320, - 64'd167011680256, 64'd6088892928, 64'd6013684224, 64'd505082688, - 64'd174943797248, - 64'd170815324160, 64'd1695074048, 64'd5749549056, 64'd598913920, - 64'd89190154240, - 64'd171721965568, - 64'd2565707008, 64'd5404309504, 64'd679595200, - 64'd3691991296, - 64'd169810132992, - 64'd6630496768, 64'd4986481152, 64'd746391296, 64'd80169967616, - 64'd165200642048, - 64'd10441671680, 64'd4505391104, 64'd798807168, 64'd161085259776, - 64'd158053154816, - 64'd13947649024, 64'd3971005440, 64'd836586944, 64'd237832192000, - 64'd148562329600, - 64'd17103477760, 64'd3393752832, 64'd859709248, 64'd309294268416, - 64'd136953618432, - 64'd19871305728, 64'd2784346368, 64'd868379008, 64'd374474440704, - 64'd123478548480, - 64'd22220722176, 64'd2153606912, 64'd863016384, 64'd432506929152, - 64'd108409978880, - 64'd24128972800, 64'd1512292864, 64'd844242304, 64'd482666741760, - 64'd92037005312, - 64'd25581041664, 64'd870935104, 64'd812862080, 64'd524376375296, - 64'd74659897344, - 64'd26569621504, 64'd239681664, 64'd769845952, 64'd557210140672, - 64'd56584978432, - 64'd27094951936, - 64'd371845536, 64'd716308672, 64'd580896161792, - 64'd38119600128, - 64'd27164561408, - 64'd954681536, 64'd653486912, 64'd595315195904, - 64'd19567282176, - 64'd26792882176, - 64'd1500634240, 64'd582715968, 64'd600498044928, - 64'd1223063168, - 64'd26000803840, - 64'd2002384256, 64'd505405504, 64'd596619952128, 64'd16630842368, - 64'd24815104000, - 64'd2453567488, 64'd423015232, 64'd583993196544, 64'd33729054720, - 64'd23267842048, - 64'd2848840704, 64'd337030624, 64'd563057786880, 64'd49826627584, - 64'd21395662848, - 64'd3183928064, 64'd248938832, 64'd534370353152, 64'd64702210048, - 64'd19239073792, - 64'd3455651072, 64'd160205840, 64'd498591858688, 64'd78160740352, - 64'd16841673728, - 64'd3661937664, 64'd72254360, 64'd456473706496, 64'd90035634176, - 64'd14249368576, - 64'd3801817344, - 64'd13556562, 64'd408843091968, 64'd100190420992, - 64'd11509573632, - 64'd3875396352, - 64'd95950400, 64'd356587700224, 64'd108519923712, - 64'd8670417920, - 64'd3883819008, - 64'd173750016, 64'd300639846400, 64'd114950856704, - 64'd5779971072, - 64'd3829213440, - 64'd245892384, 64'd241960419328, 64'd119441907712, - 64'd2885491200, - 64'd3714623232, - 64'd311441088, 64'd181523120128, 64'd121983336448, - 64'd32715716, - 64'd3543929344, - 64'd369596384, 64'd120298782720, 64'd122596114432, 64'd2734803712, - 64'd3321759488, - 64'd419702784, 64'd59240333312, 64'd121330532352, 64'd5376306176, - 64'd3053389312, - 64'd461254144, - 64'd731416192, 64'd118264520704, 64'd7854364160, - 64'd2744639488, - 64'd493896352, - 64'd58741088256, 64'd113501454336, 64'd10135356416, - 64'd2401764352, - 64'd517427488, - 64'd113970864128, 64'd107167793152, 64'd12189862912, - 64'd2031339264, - 64'd531795584, - 64'd165671337984, 64'd99410255872, 64'd13992983552, - 64'd1640147840, - 64'd537094144, - 64'd213170946048, 64'd90392961024, 64'd15524575232, - 64'd1235068032, - 64'd533555648, - 64'd255883870208, 64'd80294240256, 64'd16769404928, - 64'd822961600, - 64'd521543200, - 64'd293316329472, 64'd69303451648, 64'd17717221376, - 64'd410567744, - 64'd501540064, - 64'd325071339520, 64'd57617629184, 64'd18362755072, - 64'd4401630, - 64'd474138144, - 64'd350851596288, 64'd45438197760, 64'd18705618944, 64'd389339424, - 64'd440024864, - 64'd370460917760, 64'd32967698432, 64'd18750169088, 64'd764861952, - 64'd399969216, - 64'd383804112896, 64'd20406595584, 64'd18505261056, 64'd1116853120, - 64'd354806880, - 64'd390884950016, 64'd7950255616, 64'd17983975424, 64'd1440547328, - 64'd305424896, - 64'd391803043840, - 64'd4213928448, 64'd17203263488, 64'd1731781888, - 64'd252746048, - 64'd386749202432, - 64'd15909174272, 64'd16183558144, 64'd1987041664, - 64'd197713280, - 64'd375999365120, - 64'd26971701248, 64'd14948338688, 64'd2203492096, - 64'd141274192, - 64'd359907786752, - 64'd37252841472, 64'd13523662848, 64'd2379000320, - 64'd84366160, - 64'd338898780160, - 64'd46620835840, 64'd11937680384, 64'd2512144384, - 64'd27902050, - 64'd313458130944, - 64'd54962319360, 64'd10220119040, 64'd2602212096, 64'd27243218, - 64'd284123299840, - 64'd62183481344, 64'd8401773568, 64'd2649188096, 64'd80245000, - 64'd251473739776, - 64'd68210851840, 64'd6513990144, 64'd2653730304, 64'd130340104, - 64'd216120344576, - 64'd72991768576, 64'd4588161536, 64'd2617136384, 64'd176836592, - 64'd178695159808, - 64'd76494503936, 64'd2655238656, 64'd2541304064, 64'd219122144, - 64'd139840864256, - 64'd78708088832, 64'd745262912, 64'd2428679424, 64'd256670928, - 64'd100200562688, - 64'd79641739264, - 64'd1113069184, 64'd2282201088, 64'd289048864, - 64'd60407840768, - 64'd79324094464, - 64'd2892806656, 64'd2105238400, 64'd315917216, - 64'd21077354496, - 64'd77802110976, - 64'd4569103872, 64'd1901523584, 64'd337034816, 64'd17204037632, - 64'd75139710976, - 64'd6119537152, 64'd1675082368, 64'd352258336, 64'd53885362176, - 64'd71416266752, - 64'd7524370432, 64'd1430161280, 64'd361541280, 64'd88458821632, - 64'd66724818944, - 64'd8766772224, 64'd1171153920, 64'd364931584, 64'd120466178048, - 64'd61170216960, - 64'd9832982528, 64'd902527872, 64'd362567392, 64'd149504163840, - 64'd54867099648, - 64'd10712419328, 64'd628753024, 64'd354672160, 64'd175228796928, - 64'd47937769472, - 64'd11397739520, 64'd354231488, 64'd341548192, 64'd197358780416, - 64'd40510091264, - 64'd11884845056, 64'd83231856, 64'd323569152, 64'd215677616128, - 64'd32715292672, - 64'd12172835840, - 64'd180172848, 64'd301172096, 64'd230034898944, - 64'd24685850624, - 64'd12263920640, - 64'd432161888, 64'd274848320, 64'd240346251264, - 64'd16553392128, - 64'd12163275776, - 64'd669217728, 64'd245134048, 64'd246592552960, - 64'd8446690816, - 64'd11878867968, - 64'd888170560, 64'd212600496, 64'd248817893376, - 64'd489775968, - 64'd11421236224, - 64'd1086235904, 64'd177843856, 64'd247126884352, 64'd7199825408, - 64'd10803245056, - 64'd1261044992, 64'd141475104, 64'd241680891904, 64'd14512684032, - 64'd10039804928, - 64'd1410667520, 64'd104110152, 64'd232693678080, 64'd21348886528, - 64'd9147576320, - 64'd1533627520, 64'd66359960, 64'd220426354688, 64'd27619258368, - 64'd8144650752, - 64'd1628909952, 64'd28821298, 64'd205181698048, 64'd33246382080, - 64'd7050222080, - 64'd1695962624, - 64'd7932100, 64'd187298070528, 64'd38165393408, - 64'd5884255744, - 64'd1734687744, - 64'd43357656, 64'd167143030784, 64'd42324561920, - 64'd4667152384, - 64'd1745429632, - 64'd76951352, 64'd145106616320, 64'd45685649408, - 64'd3419417088, - 64'd1728953472, - 64'd108254256, 64'd121594593280, 64'd48224038912, - 64'd2161339904, - 64'd1686420352, - 64'd136858144, 64'd97021640704, 64'd49928663040, - 64'd912688192, - 64'd1619355392, - 64'd162410176, 64'd71804624896, 64'd50801717248, 64'd307581728, - 64'd1529612416, - 64'd184616448, 64'd46356127744, 64'd50858168320, 64'd1481589760, - 64'd1419333760, - 64'd203244672, 64'd21078155264, 64'd50125090816, 64'd2592772864, - 64'd1290908032, - 64'd218125648, - 64'd3643667456, 64'd48640860160, 64'd3626097664, - 64'd1146924288, - 64'd229153872, - 64'd27445524480, 64'd46454153216, 64'd4568240128, - 64'd990125760, - 64'd236286912, - 64'd49990291456, 64'd43622846464, 64'd5407735808, - 64'd823361984, - 64'd239544096, - 64'd70971834368, 64'd40212836352, 64'd6135093248, - 64'd649540928, - 64'd239004064, - 64'd90118692864, 64'd36296716288, 64'd6742875648, - 64'd471582400, - 64'd234801584, - 64'd107197112320, 64'd31952439296, 64'd7225745408, - 64'd292372320, - 64'd227123632, - 64'd122013368320, 64'd27261941760, 64'd7580477440, - 64'd114718976, - 64'd216204656, - 64'd134415384576, 64'd22309724160, 64'd7805936128, 64'd58687512, - 64'd202321472, - 64'd144293707776, 64'd17181462528, 64'd7903024128, 64'd225313088, - 64'd185787472, - 64'd151581720576, 64'd11962642432, 64'd7874598400, 64'd382813664, - 64'd166946560, - 64'd156255223808, 64'd6737245696, 64'd7725361664, 64'd529064992, - 64'd146166848, - 64'd158331387904, 64'd1586496384, 64'd7461724672, 64'd662188224, - 64'd123834096, - 64'd157867048960, - 64'd3412300288, 64'd7091653120, 64'd780570624, - 64'd100345176, - 64'd154956480512, - 64'd8186822656, 64'd6624487424, 64'd882881728, - 64'd76101528, - 64'd149728690176, - 64'd12670684160, 64'd6070755840, 64'd968084352, - 64'd51502828, - 64'd142344208384, - 64'd16804258816, 64'd5441968640, 64'd1035440832, - 64'd26940826, - 64'd132991549440, - 64'd20535373824, 64'd4750409216, 64'd1084514176, - 64'd2793569, - 64'd121883320320, - 64'd23819872256, 64'd4008914176, 64'd1115165056, 64'd20580006, - 64'd109252124672, - 64'd26622011392, 64'd3230659840, 64'd1127543552, 64'd42844976, - 64'd95346270208, - 64'd28914745344, 64'd2428945152, 64'd1122077440, 64'd63694820, - 64'd80425385984, - 64'd30679842816, 64'd1616980608, 64'd1099455744, 64'd82855200, - 64'd64756006912, - 64'd31907868672, 64'd807688704, 64'd1060610112, 64'd100087128, - 64'd48607227904, - 64'd32598034432, 64'd13512165, 64'd1006691072, 64'd115189488, - 64'd32246421504, - 64'd32757919744, - 64'd753761856, 64'd939043776, 64'd128000856, - 64'd15935166464, - 64'd32403066880, - 64'd1483162240, 64'd859180288, 64'd138400672, 64'd74618512, - 64'd31556468736, - 64'd2164676096, 64'd768750464, 64'd146309760, 64'd15544250368, - 64'd30247966720, - 64'd2789371904, 64'd669511808, 64'd151690080, 64'd30251536384, - 64'd28513552384, - 64'd3349500416, 64'd563298944, 64'd154544048, 64'd43993653248, - 64'd26394601472, - 64'd3838575360, 64'd451992000, 64'd154913040, 64'd56589647872, - 64'd23937046528, - 64'd4251430912, 64'd337486560, 64'd152875456, 64'd67882487808, - 64'd21190518784, - 64'd4584256512, 64'd221663488, 64'd148544336, 64'd77740703744, - 64'd18207447040, - 64'd4834612224, 64'd106360376, 64'd142064320, 64'd86059532288, - 64'd15042149376, - 64'd5001415680, - 64'd6655432, 64'd133608432, 64'd92761669632, - 64'd11749935104, - 64'd5084918784, - 64'd115711832, 64'd123374440, 64'd97797521408, - 64'd8386205184, - 64'd5086653952, - 64'd219254640, 64'd111580928, 64'd101145042944, - 64'd5005594624, - 64'd5009368576, - 64'd315867680, 64'd98463200, 64'd102809133056, - 64'd1661150336, - 64'd4856942592, - 64'd404289984, 64'd84269136, 64'd102820667392, 64'd1596436608, - 64'd4634288128, - 64'd483430176, 64'd69254864, 64'd101235122176, 64'd4719538176, - 64'd4347238912, - 64'd552377600, 64'd53680552, 64'd98130878464, 64'd7664223744, - 64'd4002430464, - 64'd610410112, 64'd37806244, 64'd93607264256, 64'd10390815744, - 64'd3607167488, - 64'd656999424, 64'd21887816, 64'd87782260736, 64'd12864362496, - 64'd3169290496, - 64'd691811968, 64'd6173181, 64'd80790077440, 64'd15055016960, - 64'd2697033984, - 64'd714708224, - 64'd9101296, 64'd72778498048, 64'd16938331136, - 64'd2198887424, - 64'd725737856, - 64'd23714064, 64'd63906152448, 64'd18495447040, - 64'd1683453824, - 64'd725132608, - 64'd37461312, 64'd54339653632, 64'd19713210368, - 64'd1159312768, - 64'd713296768, - 64'd50159536, 64'd44250787840, 64'd20584165376, - 64'd634889024, - 64'd690794752, - 64'd61647676, 64'd33813639168, 64'd21106491392, - 64'd118326248, - 64'd658337280, - 64'd71788872, 64'd23201835008, 64'd21283842048, 64'd382629120, - 64'd616765184, - 64'd80471752, 64'd12585860096, 64'd21125087232, 64'd860734720, - 64'd567032064, - 64'd87611304, 64'd2130512896, 64'd20644018176, 64'd1309347456, - 64'd510185696, - 64'd93149288, - 64'd8007448576, 64'd19858956288, 64'd1722505984, - 64'd447348576, - 64'd97054256, - 64'd17681471488, 64'd18792316928, 64'd2095000448, - 64'd379698048, - 64'd99321104, - 64'd26757134336, 64'd17470130176, 64'd2422427648, - 64'd308446240, - 64'd99970280, - 64'd35113828352, 64'd15921509376, 64'd2701231360, - 64'd234820016, - 64'd99046608, - 64'd42646147072, 64'd14178094080, 64'd2928730368, - 64'd160041504, - 64'd96617760, - 64'd49265025024, 64'd12273478656, 64'd3103128832, - 64'd85309368, - 64'd92772416, - 64'd54898561024, 64'd10242625536, 64'd3223515136, - 64'd11780941, - 64'd87618232, - 64'd59492548608, 64'd8121272832, 64'd3289845760, 64'd59444232, - 64'd81279464, - 64'd63010721792, 64'd5945358336, 64'd3302916864, 64'd127339528, - 64'd73894544, - 64'd65434730496, 64'd3750452736, 64'd3264323072, 64'd190964656, - 64'd65613412, - 64'd66763780096, 64'd1571222144, 64'd3176407040, 64'd249477360, - 64'd56594828, - 64'd67014103040, - 64'd559078976, 64'd3042195712, 64'd302143104, - 64'd47003604, - 64'd66218090496, - 64'd2609076224, 64'd2865332736, 64'd348342816, - 64'd37007848, - 64'd64423264256, - 64'd4549698048, 64'd2649999360, 64'd387578592, - 64'd26776244, - 64'd61691031552, - 64'd6354548224, 64'd2400832000, 64'd419477408, - 64'd16475429, - 64'd58095259648, - 64'd8000225280, 64'd2122835328, 64'd443792480, - 64'd6267468, - 64'd53720711168, - 64'd9466584064, 64'd1821291904, 64'd460403008, 64'd3692493, - 64'd48661364736, - 64'd10736937984, 64'd1501670912, 64'd469311648, 64'd13258402, - 64'd43018645504, - 64'd11798201344, 64'd1169537280, 64'd470640448, 64'd22295256, - 64'd36899602432, - 64'd12640969728, 64'd830462080, 64'd464624800, 64'd30680818, - 64'd30415069184, - 64'd13259542528, 64'd489935872, 64'd451606016, 64'd38307084, - 64'd23677794304, - 64'd13651887104, 64'd153286496, 64'd432022368, 64'd45081468, - 64'd16800658432, - 64'd13819544576, - 64'd174398144, 64'd406399232, 64'd50927724, - 64'd9894899712, - 64'd13767486464, - 64'd488340800, 64'd375337760, 64'd55786572, - 64'd3068452864, - 64'd13503922176, - 64'd784138432, 64'd339503104, 64'd59616036, 64'd3575611392, - 64'd13040061440, - 64'd1057817792, 64'd299612032, 64'd62391524, 64'd9940521984, - 64'd12389841920, - 64'd1305882624, 64'd256419936, 64'd64105612, 64'd15937092608, - 64'd11569616896, - 64'd1525351552, 64'd210707840, 64'd64767576, 64'd21484853248, - 64'd10597824512, - 64'd1713787136, 64'd163269520, 64'd64402692, 64'd26512994304, - 64'd9494629376, - 64'd1869315200, 64'd114898680, 64'd63051300, 64'd30961149952, - 64'd8281552384, - 64'd1990634752, 64'd66376692, 64'd60767672, 64'd34779967488, - 64'd6981092352, - 64'd2077019008, 64'd18460890, 64'd57618692, 64'd37931511808, - 64'd5616342528, - 64'd2128306816, - 64'd28126356, 64'd53682408, 64'd40389468160, - 64'd4210614016, - 64'd2144887040, - 64'd72707656, 64'd49046428, 64'd42139148288, - 64'd2787066880, - 64'd2127672832, - 64'd114659568, 64'd43806252, 64'd43177336832, - 64'd1368355968, - 64'd2078070528, - 64'd153420464, 64'd38063520, 64'd43511943168, 64'd23702650, - 64'd1997940864, - 64'd188497136, 64'd31924228, 64'd43161522176, 64'd1368441600, - 64'd1889554944, - 64'd219470112, 64'd25496940, 64'd42154598400, 64'd2646623744, - 64'd1755545344, - 64'd245997696, 64'd18891022, 64'd40528924672, 64'd3840692224, - 64'd1598852736, - 64'd267818624, 64'd12214913, 64'd38330544128, 64'd4934985728, - 64'd1422670208, - 64'd284753408, 64'd5574480, 64'd35612844032, 64'd5915916800, - 64'd1230385152, - 64'd296704352, - 64'd928537, 64'd32435431424, 64'd6772112896, - 64'd1025520192, - 64'd303654304, - 64'd7197964, 64'd28863043584, 64'd7494518784, - 64'd811674048, - 64'd305664192, - 64'd13144493, 64'd24964341760, 64'd8076455424, - 64'd592463360, - 64'd302869440, - 64'd18686836, 64'd20810729472, 64'd8513648640, - 64'd371465760, - 64'd295475424, - 64'd23752716, 64'd16475149312, 64'd8804207616, - 64'd152165872, - 64'd283751840, - 64'd28279676, 64'd12030904320, 64'd8948580352, 64'd62095476, - 64'd268026352, - 64'd32215728, 64'd7550502912, 64'd8949464064, 64'd268168304, - 64'd248677680, - 64'd35519788, 64'd3104569856, 64'd8811685888, 64'd463135744, - 64'd226127840, - 64'd38161968, - 64'd1239189120, 64'd8542060544, 64'd644351488, - 64'd200834240, - 64'd40123628, - 64'd5416935936, 64'd8149216256, 64'd809471616, - 64'd173281424, - 64'd41397324, - 64'd9369559040, 64'd7643397120, 64'd956480640, - 64'd143972544, - 64'd41986520, - 64'd13043429376, 64'd7036254208, 64'd1083711744, - 64'd113421008, - 64'd41905164, - 64'd16391049216, 64'd6340613120, 64'd1189860736, - 64'd82142176, - 64'd41177136, - 64'd19371575296, 64'd5570238976, 64'd1273994496, - 64'd50645276, - 64'd39835528, - 64'd21951229952, 64'd4739590656, 64'd1335551872, - 64'd19425748, - 64'd37921832, - 64'd24103593984, 64'd3863571968, 64'd1374341120, 64'd11041996, - 64'd35484996, - 64'd25809750016, 64'd2957286656, 64'd1390529536, 64'd40311192, - 64'd32580432, - 64'd27058341888, 64'd2035798272, 64'd1384628608, 64'd67968728, - 64'd29268928, - 64'd27845476352, 64'd1113897088, 64'd1357475456, 64'd93640400, - 64'd25615532, - 64'd28174551040, 64'd205880560, 64'd1310208000, 64'd116995408, - 64'd21688388, - 64'd28055937024, - 64'd674651648, 64'd1244237184, 64'd137750016, - 64'd17557590, - 64'd27506599936, - 64'd1514984704, 64'd1161216512, 64'd155670336, - 64'd13294021, - 64'd26549600256, - 64'd2303456000, 64'd1063007808, 64'd170574336, - 64'd8968230, - 64'd25213538304, - 64'd3029600256, 64'd951645312, 64'd182332832, - 64'd4649348, - 64'd23531919360, - 64'd3684270848, 64'd829298368, 64'd190869744, - 64'd404071, - 64'd21542475776, - 64'd4259737856, 64'd698233472, 64'd196161488, 64'd3704301, - 64'd19286431744, - 64'd4749759488, 64'd560775680, 64'd198235584, 64'd7616722, - 64'd16807752704, - 64'd5149628416, 64'd419270496, 64'd197168432, 64'd11279177, - 64'd14152366080, - 64'd5456193024, 64'd276047136, 64'd193082576, 64'd14643346, - 64'd11367388160, - 64'd5667854336, 64'd133382744, 64'd186143184, 64'd17667162, - 64'd8500353536, - 64'd5784537600, - 64'd6531030, 64'd176554064, 64'd20315252, - 64'd5598459904, - 64'd5807642112, - 64'd141619152, 64'd164553216, 64'd22559258, - 64'd2707853312, - 64'd5739970048, - 64'd269951392, 64'd150407984, 64'd24378042, 64'd127054280, - 64'd5585635840, - 64'd389767392, 64'd134409888, 64'd25757768, 64'd2864213504, - 64'd5349958144, - 64'd499498080, 64'd116869344, 64'd26691872, 64'd5464509952, - 64'd5039334912, - 64'd597783744, 64'd98110200, 64'd27180914};
endpackage
`endif
