`ifndef COEFFICIENTS_FX_SV_
`define COEFFICIENTS_FX_SV_
package Coefficients_Fx;
	localparam N = 4;
	localparam M = 4;
	localparam COEFF_BIAS = 48;
	localparam logic signed[63:0] Lfr[0:3] = {64'd278939910093526, 64'd278939910093526, 64'd275816626731508, 64'd275816626731508};
	localparam logic signed[63:0] Lfi[0:3] = {64'd11276861423257, - 64'd11276861423257, 64'd4532123198530, - 64'd4532123198530};
	localparam logic signed[63:0] Lbr[0:3] = {64'd278939910093526, 64'd278939910093526, 64'd275816626731508, 64'd275816626731508};
	localparam logic signed[63:0] Lbi[0:3] = {64'd11276861423257, - 64'd11276861423257, 64'd4532123198530, - 64'd4532123198530};
	localparam logic signed[63:0] Wfr[0:3] = {- 64'd1795674633, - 64'd1795674633, - 64'd533851843, - 64'd533851843};
	localparam logic signed[63:0] Wfi[0:3] = {- 64'd70718785, 64'd70718785, - 64'd1029591743, 64'd1029591743};
	localparam logic signed[63:0] Wbr[0:3] = {64'd1795674633, 64'd1795674633, 64'd533851843, 64'd533851843};
	localparam logic signed[63:0] Wbi[0:3] = {64'd70718785, - 64'd70718785, 64'd1029591743, - 64'd1029591743};
	localparam logic signed[63:0] Ffr[0:3][0:99] = '{
		'{- 64'd88776608138663776, - 64'd7242245853080698, 64'd673217222953428, - 64'd5885714537304, - 64'd92292018980244400, - 64'd6818568896873604, 64'd676486126205592, - 64'd7478244584595, - 64'd95594412957760064, - 64'd6390311678074589, 64'd678560971769394, - 64'd9032164350417, - 64'd98681699417100496, - 64'd5958271101876197, 64'd679457755875843, - 64'd10545483994509, - 64'd101552184550611792, - 64'd5523237442249447, 64'd679194200034766, - 64'd12016314623546, - 64'd104204567774058880, - 64'd5085993117652344, 64'd677789692985040, - 64'd13442869828075, - 64'd106637937499688576, - 64'd4647311499972762, 64'd675265230781322, - 64'd14823467021539, - 64'd108851766322379328, - 64'd4207955758171454, 64'd671643355148691, - 64'd16156528582381, - 64'd110845905636577824, - 64'd3768677738008483, 64'd666948090237456, - 64'd17440582800506, - 64'd112620579702391936, - 64'd3330216879152979, 64'd661204877910872, - 64'd18674264629703, - 64'd114176379179839824, - 64'd2893299170891838, 64'd654440511698840, - 64'd19856316247935, - 64'd115514254150840064, - 64'd2458636147568046, 64'd646683069550753, - 64'd20985587427663, - 64'd116635506649073344, - 64'd2026923924793884, 64'd637961845520457, - 64'd22061035718717, - 64'd117541782718345920, - 64'd1598842277398421, 64'd628307280515980, - 64'd23081726446436, - 64'd118235064020544288, - 64'd1175053759982688, 64'd617750892246058, - 64'd24046832528115, - 64'd118717659014685152, - 64'd756202870869806, 64'd606325204494687, - 64'd24955634111016, - 64'd118992193728937280, - 64'd342915260151333, 64'd594063675853948, - 64'd25807518035498, - 64'd119061602147820352, 64'd64203017554733, 64'd581000628044100, - 64'd26601977126985, - 64'd118929116237073184, 64'd464566205104279, 64'd567171173948559, - 64'd27338609320798, - 64'd118598255628926768, 64'd857609499140658, 64'd552611145489763, - 64'd28017116624032, - 64'd118072816990718832, 64'd1242789660360759, 64'd537357021470127, - 64'd28637303918901, - 64'd117356863099947136, 64'd1619585577456348, 64'd521445855500345, - 64'd29199077612148, - 64'd116454711648975328, 64'd1987498784536060, 64'd504915204135132, - 64'd29702444135316, - 64'd115370923802683104, 64'd2346053931915101, 64'd487803055334201, - 64'd30147508300851, - 64'd114110292532387648, 64'd2694799210240125, 64'd470147757363787, - 64'd30534471519142},
		'{- 64'd88776608138727552, - 64'd7242245853076649, 64'd673217222953349, - 64'd5885714537298, - 64'd92292018980305536, - 64'd6818568896869722, 64'd676486126205516, - 64'd7478244584589, - 64'd95594412957818496, - 64'd6390311678070879, 64'd678560971769321, - 64'd9032164350412, - 64'd98681699417156176, - 64'd5958271101872662, 64'd679457755875774, - 64'd10545483994503, - 64'd101552184550664640, - 64'd5523237442246090, 64'd679194200034700, - 64'd12016314623541, - 64'd104204567774108896, - 64'd5085993117649168, 64'd677789692984977, - 64'd13442869828070, - 64'd106637937499735712, - 64'd4647311499969770, 64'd675265230781262, - 64'd14823467021535, - 64'd108851766322423552, - 64'd4207955758168646, 64'd671643355148634, - 64'd16156528582377, - 64'd110845905636619088, - 64'd3768677738005862, 64'd666948090237403, - 64'd17440582800501, - 64'd112620579702430256, - 64'd3330216879150546, 64'd661204877910822, - 64'd18674264629699, - 64'd114176379179875136, - 64'd2893299170889594, 64'd654440511698794, - 64'd19856316247931, - 64'd115514254150872384, - 64'd2458636147565992, 64'd646683069550711, - 64'd20985587427659, - 64'd116635506649102656, - 64'd2026923924792021, 64'd637961845520418, - 64'd22061035718713, - 64'd117541782718372256, - 64'd1598842277396749, 64'd628307280515945, - 64'd23081726446433, - 64'd118235064020567616, - 64'd1175053759981206, 64'd617750892246026, - 64'd24046832528112, - 64'd118717659014705504, - 64'd756202870868512, 64'd606325204494658, - 64'd24955634111014, - 64'd118992193728954656, - 64'd342915260150229, 64'd594063675853922, - 64'd25807518035496, - 64'd119061602147834784, 64'd64203017555650, 64'd581000628044078, - 64'd26601977126983, - 64'd118929116237084704, 64'd464566205105010, 64'd567171173948541, - 64'd27338609320796, - 64'd118598255628935360, 64'd857609499141205, 64'd552611145489749, - 64'd28017116624031, - 64'd118072816990724560, 64'd1242789660361124, 64'd537357021470116, - 64'd28637303918900, - 64'd117356863099950048, 64'd1619585577456533, 64'd521445855500337, - 64'd29199077612147, - 64'd116454711648975456, 64'd1987498784536068, 64'd504915204135127, - 64'd29702444135315, - 64'd115370923802680480, 64'd2346053931914935, 64'd487803055334200, - 64'd30147508300851, - 64'd114110292532382336, 64'd2694799210239788, 64'd470147757363789, - 64'd30534471519142},
		'{- 64'd88355216767193600, - 64'd7210717608321972, 64'd652814047329850, - 64'd74474048717025, - 64'd91858913475248672, - 64'd6806001903237092, 64'd622973704183345, - 64'd72155440125182, - 64'd95163132456448672, - 64'd6412774464623528, 64'd593900038914348, - 64'd69880647819613, - 64'd98273569487507344, - 64'd6030841880384146, 64'd565582022235033, - 64'd67649448246895, - 64'd101195823672693504, - 64'd5660010893658376, 64'd538008559703970, - 64'd65461597775446, - 64'd103935397552176256, - 64'd5300088524883438, 64'd511168501662055, - 64'd63316833651065, - 64'd106497697270143200, - 64'd4950882188845119, 64'd485050652812178, - 64'd61214874927375, - 64'd108888032800216368, - 64'd4612199806838576, 64'd459643781450378, - 64'd59155423371540, - 64'd111111618225751072, - 64'd4283849914058110, 64'd434936628356130, - 64'd57138164345637, - 64'd113173572072661216, - 64'd3965641762333352, 64'd410917915349351, - 64'd55162767664057, - 64'd115078917692473632, - 64'd3657385418327684, 64'd387576353521621, - 64'd53228888427322, - 64'd116832583693370816, - 64'd3358891857313212, 64'd364900651149051, - 64'd51336167832687, - 64'd118439404417039040, - 64'd3069973052634992, 64'd342879521294128, - 64'd49484233961915, - 64'd119904120459193856, - 64'd2790442060975596, 64'd321501689103792, - 64'd47672702546602, - 64'd121231379231710912, - 64'd2520113103529546, 64'd300755898810927, - 64'd45901177711433, - 64'd122425735564343952, - 64'd2258801643195464, 64'd280630920446329, - 64'd44169252695746, - 64'd123491652344065504, - 64'd2006324457892246, 64'd261115556268174, - 64'd42476510553788, - 64'd124433501190118432, - 64'd1762499710103830, 64'd242198646915861, - 64'd40822524834034, - 64'd125255563162918528, - 64'd1527147012755594, 64'd223869077295067, - 64'd39206860237959, - 64'd125962029504999408, - 64'd1300087491523733, 64'd206115782200739, - 64'd37629073258616, - 64'd126557002412241056, - 64'd1081143843677293, 64'd188927751684637, - 64'd36088712799422, - 64'd127044495833673088, - 64'd870140393550984, 64'd172294036173990, - 64'd34585320773506, - 64'd127428436298192192, - 64'd666903144745155, 64'd156203751347696, - 64'd33118432683989, - 64'd127712663766581200, - 64'd471259829147740, 64'd140646082776425, - 64'd31687578185584, - 64'd127900932507263808, - 64'd283039952871314, 64'd125610290332884, - 64'd30292281627854},
		'{- 64'd88355216767386768, - 64'd7210717608309690, 64'd652814047329616, - 64'd74474048717007, - 64'd91858913475437136, - 64'd6806001903225109, 64'd622973704183117, - 64'd72155440125165, - 64'd95163132456632496, - 64'd6412774464611841, 64'd593900038914125, - 64'd69880647819597, - 64'd98273569487686592, - 64'd6030841880372750, 64'd565582022234815, - 64'd67649448246879, - 64'd101195823672868208, - 64'd5660010893647267, 64'd538008559703758, - 64'd65461597775430, - 64'd103935397552346496, - 64'd5300088524872613, 64'd511168501661848, - 64'd63316833651049, - 64'd106497697270309040, - 64'd4950882188834574, 64'd485050652811977, - 64'd61214874927360, - 64'd108888032800377888, - 64'd4612199806828306, 64'd459643781450182, - 64'd59155423371526, - 64'd111111618225908304, - 64'd4283849914048112, 64'd434936628355939, - 64'd57138164345623, - 64'd113173572072814240, - 64'd3965641762323622, 64'd410917915349164, - 64'd55162767664043, - 64'd115078917692622528, - 64'd3657385418318216, 64'd387576353521439, - 64'd53228888427309, - 64'd116832583693515648, - 64'd3358891857304003, 64'd364900651148874, - 64'd51336167832674, - 64'd118439404417179840, - 64'd3069973052626038, 64'd342879521293956, - 64'd49484233961902, - 64'd119904120459330720, - 64'd2790442060966894, 64'd321501689103625, - 64'd47672702546590, - 64'd121231379231843888, - 64'd2520113103521090, 64'd300755898810764, - 64'd45901177711421, - 64'd122425735564473120, - 64'd2258801643187250, 64'd280630920446172, - 64'd44169252695734, - 64'd123491652344190928, - 64'd2006324457884270, 64'd261115556268021, - 64'd42476510553776, - 64'd124433501190240176, - 64'd1762499710096088, 64'd242198646915712, - 64'd40822524834023, - 64'd125255563163036640, - 64'd1527147012748084, 64'd223869077294923, - 64'd39206860237948, - 64'd125962029505113984, - 64'd1300087491516448, 64'd206115782200599, - 64'd37629073258605, - 64'd126557002412352128, - 64'd1081143843670230, 64'd188927751684501, - 64'd36088712799412, - 64'd127044495833780736, - 64'd870140393544138, 64'd172294036173858, - 64'd34585320773496, - 64'd127428436298296480, - 64'd666903144738522, 64'd156203751347568, - 64'd33118432683980, - 64'd127712663766682176, - 64'd471259829141318, 64'd140646082776301, - 64'd31687578185574, - 64'd127900932507361568, - 64'd283039952865098, 64'd125610290332764, - 64'd30292281627845}};
	localparam logic signed[63:0] Ffi[0:3][0:99] = '{
		'{64'd107703265549738064, - 64'd8947071520977922, - 64'd232934047530405, 64'd41073311006417, 64'd103176552463027872, - 64'd9156640347428454, - 64'd203864747109806, 64'd40467587652981, 64'd98549769089416768, - 64'd9347347755640880, - 64'd174926291869582, 64'd39803517402087, 64'd93832350891096016, - 64'd9519180117281880, - 64'd146165341452405, 64'd39083172608701, 64'd89033732109869584, - 64'd9672155853539060, - 64'd117627494402776, 64'd38308686683285, 64'd84163329879103072, - 64'd9806324880801568, - 64'd89357228603024, 64'd37482249497631, 64'd79230528623918016, - 64'd9921768012283748, - 64'd61397844571438, 64'd36606102770485, 64'd74244664771229408, - 64'd10018596317320144, - 64'd33791411671403, 64'd35682535441095, 64'd69215011790349648, - 64'd10096950440103238, - 64'd6578717274732, 64'd34713879038661, 64'd64150765583986400, - 64'd10156999879674868, 64'd20200781083337, 64'd33702503055577, 64'd59061030248547488, - 64'd10198942233017976, 64'd46509000525631, 64'd32650810332197, 64'd53954804221733768, - 64'd10223002403127416, 64'd72309274604807, 64'd31561232460715, 64'd48840966834455424, - 64'd10229431773966964, 64'd97566392004763, 64'd30436225215614, 64'd43728265283145904, - 64'd10218507354244318, 64'd122246632156539, 64'd29278264017934, 64'd38625302037577456, - 64'd10190530891956972, 64'd146317797759052, 64'd28089839440465, 64'd33540522698301016, - 64'd10145827961679208, 64'd169749244200350, 64'd26873452760785, 64'd28482204316844112, - 64'd10084747026574258, 64'd192511905880381, 64'd25631611568843, 64'd23458444190805936, - 64'd10007658477125936, 64'd214578319441481, 64'd24366825435609, 64'd18477149144990256, - 64'd9914953648590698, 64'd235922643917893, 64'd23081601649110, 64'd13546025308714328, - 64'd9807043819174324, 64'd256520677820646, 64'd21778441023919, 64'd8672568398431088, - 64'd9684359190937200, 64'd276349873179018, 64'd20459833789988, 64'd3864054513799336, - 64'd9547347855428568, 64'd295389346564595, 64'd19128255566438, - 64'd872468545660632, - 64'd9396474746043208, 64'd313619887128605, 64'd17786163425729, - 64'd5530189437183984, - 64'd9232220579083878, 64'd331023961687728, 64'd16435992053359, - 64'd10102540899496720, - 64'd9055080785499432, 64'd347585716898006, 64'd15080150008005},
		'{- 64'd107703265549686464, 64'd8947071520974648, 64'd232934047530462, - 64'd41073311006421, - 64'd103176552462974192, 64'd9156640347425048, 64'd203864747109865, - 64'd40467587652985, - 64'd98549769089361104, 64'd9347347755637348, 64'd174926291869644, - 64'd39803517402091, - 64'd93832350891038528, 64'd9519180117278230, 64'd146165341452470, - 64'd39083172608705, - 64'd89033732109810368, 64'd9672155853535304, 64'd117627494402843, - 64'd38308686683290, - 64'd84163329879042272, 64'd9806324880797710, 64'd89357228603093, - 64'd37482249497635, - 64'd79230528623855760, 64'd9921768012279798, 64'd61397844571508, - 64'd36606102770490, - 64'd74244664771165840, 64'd10018596317316110, 64'd33791411671475, - 64'd35682535441100, - 64'd69215011790284872, 64'd10096950440099126, 64'd6578717274805, - 64'd34713879038666, - 64'd64150765583920560, 64'd10156999879670690, - 64'd20200781083262, - 64'd33702503055583, - 64'd59061030248480696, 64'd10198942233013736, - 64'd46509000525554, - 64'd32650810332202, - 64'd53954804221666176, 64'd10223002403123124, - 64'd72309274604729, - 64'd31561232460721, - 64'd48840966834387152, 64'd10229431773962628, - 64'd97566392004684, - 64'd30436225215620, - 64'd43728265283077064, 64'd10218507354239948, - 64'd122246632156459, - 64'd29278264017939, - 64'd38625302037508176, 64'd10190530891952574, - 64'd146317797758972, - 64'd28089839440471, - 64'd33540522698231432, 64'd10145827961674790, - 64'd169749244200269, - 64'd26873452760791, - 64'd28482204316774328, 64'd10084747026569828, - 64'd192511905880300, - 64'd25631611568849, - 64'd23458444190736088, 64'd10007658477121504, - 64'd214578319441399, - 64'd24366825435615, - 64'd18477149144920448, 64'd9914953648586268, - 64'd235922643917811, - 64'd23081601649116, - 64'd13546025308644696, 64'd9807043819169904, - 64'd256520677820564, - 64'd21778441023925, - 64'd8672568398361736, 64'd9684359190932798, - 64'd276349873178936, - 64'd20459833789994, - 64'd3864054513730376, 64'd9547347855424192, - 64'd295389346564514, - 64'd19128255566444, 64'd872468545729080, 64'd9396474746038864, - 64'd313619887128524, - 64'd17786163425735, 64'd5530189437251816, 64'd9232220579079572, - 64'd331023961687648, - 64'd16435992053364, 64'd10102540899563848, 64'd9055080785495172, - 64'd347585716897926, - 64'd15080150008011},
		'{64'd327914229854852992, - 64'd16132963874025046, 64'd1038246167410144, - 64'd51020251934053, 64'd319899697871776704, - 64'd15924753197771214, 64'd1027886004934731, - 64'd51193749141451, 64'd311989863798591104, - 64'd15714211612504252, 64'd1017253638204449, - 64'd51326425925515, 64'd304185834803758720, - 64'd15501570951755914, 64'd1006366883742788, - 64'd51419808379449, 64'd296488604089275968, - 64'd15287055274431814, 64'd995243022330351, - 64'd51475388318663, 64'd288899054738239104, - 64'd15070881023600346, 64'd983898808725565, - 64'd51494623646558, 64'd281417963483320224, - 64'd14853257184054888, 64'd972350481349960, - 64'd51478938728343, 64'd274046004396780480, - 64'd14634385438593302, 64'd960613771932999, - 64'd51429724772316, 64'd266783752502675136, - 64'd14414460322961760, 64'd948703915111656, - 64'd51348340218067, 64'd259631687311931712, - 64'd14193669379412916, 64'd936635657980159, - 64'd51236111131066, 64'd252590196281004288, - 64'd13972193308831394, 64'd924423269585548, - 64'd51094331603127, 64'd245659578194833664, - 64'd13750206121382268, 64'd912080550364871, - 64'd50924264158244, 64'd238840046474860192, - 64'd13527875285641054, 64'd899620841520088, - 64'd50727140163322, 64'd232131732412860224, - 64'd13305361876166310, 64'd887057034326906, - 64'd50504160243335, 64'd225534688331392544, - 64'd13082820719478520, 64'd874401579373997, - 64'd50256494700464, 64'd219048890671661408, - 64'd12860400538411460, 64'd861666495729220, - 64'd49985283936770, 64'd212674243009616960, - 64'd12638244094804652, 64'd848863380029643, - 64'd49691638879994, 64'd206410579001130624, - 64'd12416488330507796, 64'd836003415492366, - 64'd49376641412073, 64'd200257665257095456, - 64'd12195264506670468, 64'd823097380843278, - 64'd49041344799975, 64'd194215204149316032, - 64'd11974698341292420, 64'd810155659161094, - 64'd48686774128483, 64'd188282836548062176, - 64'd11754910145012030, 64'd797188246634127, - 64'd48313926734564, 64'd182460144492173664, - 64'd11536014955112534, 64'd784204761227466, - 64'd47923772642960, 64'd176746653792611072, - 64'd11318122667727552, 64'd771214451258330, - 64'd47517255002685, 64'd171141836570357568, - 64'd11101338168229462, 64'd758226203877556, - 64'd47095290524082, 64'd165645113729583616, - 64'd10885761459785948, 64'd745248553455290, - 64'd46658769916138},
		'{- 64'd327914229854801664, 64'd16132963874021790, - 64'd1038246167410088, 64'd51020251934049, - 64'd319899697871723264, 64'd15924753197767824, - 64'd1027886004934672, 64'd51193749141447, - 64'd311989863798535680, 64'd15714211612500738, - 64'd1017253638204388, 64'd51326425925511, - 64'd304185834803701504, 64'd15501570951752284, - 64'd1006366883742724, 64'd51419808379444, - 64'd296488604089217024, 64'd15287055274428074, - 64'd995243022330285, 64'd51475388318658, - 64'd288899054738178496, 64'd15070881023596500, - 64'd983898808725497, 64'd51494623646554, - 64'd281417963483258144, 64'd14853257184050946, - 64'd972350481349890, 64'd51478938728339, - 64'd274046004396716960, 64'd14634385438589270, - 64'd960613771932928, 64'd51429724772311, - 64'd266783752502610304, 64'd14414460322957642, - 64'd948703915111582, 64'd51348340218062, - 64'd259631687311865600, 64'd14193669379408722, - 64'd936635657980084, 64'd51236111131060, - 64'd252590196280937088, 64'd13972193308827128, - 64'd924423269585471, 64'd51094331603121, - 64'd245659578194765408, 64'd13750206121377934, - 64'd912080550364793, 64'd50924264158238, - 64'd238840046474790976, 64'd13527875285636658, - 64'd899620841520008, 64'd50727140163316, - 64'd232131732412790144, 64'd13305361876161860, - 64'd887057034326825, 64'd50504160243330, - 64'd225534688331321664, 64'd13082820719474018, - 64'd874401579373915, 64'd50256494700458, - 64'd219048890671589760, 64'd12860400538406916, - 64'd861666495729137, 64'd49985283936764, - 64'd212674243009544736, 64'd12638244094800064, - 64'd848863380029560, 64'd49691638879988, - 64'd206410579001057824, 64'd12416488330503172, - 64'd836003415492282, 64'd49376641412067, - 64'd200257665257022144, 64'd12195264506665812, - 64'd823097380843194, 64'd49041344799968, - 64'd194215204149242304, 64'd11974698341287738, - 64'd810155659161008, 64'd48686774128477, - 64'd188282836547988064, 64'd11754910145007324, - 64'd797188246634041, 64'd48313926734557, - 64'd182460144492099264, 64'd11536014955107808, - 64'd784204761227379, 64'd47923772642954, - 64'd176746653792536448, 64'd11318122667722810, - 64'd771214451258244, 64'd47517255002679, - 64'd171141836570282784, 64'd11101338168224710, - 64'd758226203877469, 64'd47095290524076, - 64'd165645113729508704, 64'd10885761459781186, - 64'd745248553455202, 64'd46658769916132}};
	localparam logic signed[63:0] Fbr[0:3][0:99] = '{
		'{64'd88776608138663776, - 64'd7242245853080698, - 64'd673217222953428, - 64'd5885714537304, 64'd92292018980244400, - 64'd6818568896873604, - 64'd676486126205592, - 64'd7478244584595, 64'd95594412957760064, - 64'd6390311678074589, - 64'd678560971769394, - 64'd9032164350417, 64'd98681699417100496, - 64'd5958271101876197, - 64'd679457755875843, - 64'd10545483994509, 64'd101552184550611792, - 64'd5523237442249447, - 64'd679194200034766, - 64'd12016314623546, 64'd104204567774058880, - 64'd5085993117652344, - 64'd677789692985040, - 64'd13442869828075, 64'd106637937499688576, - 64'd4647311499972762, - 64'd675265230781322, - 64'd14823467021539, 64'd108851766322379328, - 64'd4207955758171454, - 64'd671643355148691, - 64'd16156528582381, 64'd110845905636577824, - 64'd3768677738008483, - 64'd666948090237456, - 64'd17440582800506, 64'd112620579702391936, - 64'd3330216879152979, - 64'd661204877910872, - 64'd18674264629703, 64'd114176379179839824, - 64'd2893299170891838, - 64'd654440511698840, - 64'd19856316247935, 64'd115514254150840064, - 64'd2458636147568046, - 64'd646683069550753, - 64'd20985587427663, 64'd116635506649073344, - 64'd2026923924793884, - 64'd637961845520457, - 64'd22061035718717, 64'd117541782718345920, - 64'd1598842277398421, - 64'd628307280515980, - 64'd23081726446436, 64'd118235064020544288, - 64'd1175053759982688, - 64'd617750892246058, - 64'd24046832528115, 64'd118717659014685152, - 64'd756202870869806, - 64'd606325204494687, - 64'd24955634111016, 64'd118992193728937280, - 64'd342915260151333, - 64'd594063675853948, - 64'd25807518035498, 64'd119061602147820352, 64'd64203017554733, - 64'd581000628044100, - 64'd26601977126985, 64'd118929116237073184, 64'd464566205104279, - 64'd567171173948559, - 64'd27338609320798, 64'd118598255628926768, 64'd857609499140658, - 64'd552611145489763, - 64'd28017116624032, 64'd118072816990718832, 64'd1242789660360759, - 64'd537357021470127, - 64'd28637303918901, 64'd117356863099947136, 64'd1619585577456348, - 64'd521445855500345, - 64'd29199077612148, 64'd116454711648975328, 64'd1987498784536060, - 64'd504915204135132, - 64'd29702444135316, 64'd115370923802683104, 64'd2346053931915101, - 64'd487803055334201, - 64'd30147508300851, 64'd114110292532387648, 64'd2694799210240125, - 64'd470147757363787, - 64'd30534471519142},
		'{64'd88776608138727552, - 64'd7242245853076649, - 64'd673217222953349, - 64'd5885714537298, 64'd92292018980305536, - 64'd6818568896869722, - 64'd676486126205516, - 64'd7478244584589, 64'd95594412957818496, - 64'd6390311678070879, - 64'd678560971769321, - 64'd9032164350412, 64'd98681699417156176, - 64'd5958271101872662, - 64'd679457755875774, - 64'd10545483994503, 64'd101552184550664640, - 64'd5523237442246090, - 64'd679194200034700, - 64'd12016314623541, 64'd104204567774108896, - 64'd5085993117649168, - 64'd677789692984977, - 64'd13442869828070, 64'd106637937499735712, - 64'd4647311499969770, - 64'd675265230781262, - 64'd14823467021535, 64'd108851766322423552, - 64'd4207955758168646, - 64'd671643355148634, - 64'd16156528582377, 64'd110845905636619088, - 64'd3768677738005862, - 64'd666948090237403, - 64'd17440582800501, 64'd112620579702430256, - 64'd3330216879150546, - 64'd661204877910822, - 64'd18674264629699, 64'd114176379179875136, - 64'd2893299170889594, - 64'd654440511698794, - 64'd19856316247931, 64'd115514254150872384, - 64'd2458636147565992, - 64'd646683069550711, - 64'd20985587427659, 64'd116635506649102656, - 64'd2026923924792021, - 64'd637961845520418, - 64'd22061035718713, 64'd117541782718372256, - 64'd1598842277396749, - 64'd628307280515945, - 64'd23081726446433, 64'd118235064020567616, - 64'd1175053759981206, - 64'd617750892246026, - 64'd24046832528112, 64'd118717659014705504, - 64'd756202870868512, - 64'd606325204494658, - 64'd24955634111014, 64'd118992193728954656, - 64'd342915260150229, - 64'd594063675853922, - 64'd25807518035496, 64'd119061602147834784, 64'd64203017555650, - 64'd581000628044078, - 64'd26601977126983, 64'd118929116237084704, 64'd464566205105010, - 64'd567171173948541, - 64'd27338609320796, 64'd118598255628935360, 64'd857609499141205, - 64'd552611145489749, - 64'd28017116624031, 64'd118072816990724560, 64'd1242789660361124, - 64'd537357021470116, - 64'd28637303918900, 64'd117356863099950048, 64'd1619585577456533, - 64'd521445855500337, - 64'd29199077612147, 64'd116454711648975456, 64'd1987498784536068, - 64'd504915204135127, - 64'd29702444135315, 64'd115370923802680480, 64'd2346053931914935, - 64'd487803055334200, - 64'd30147508300851, 64'd114110292532382336, 64'd2694799210239788, - 64'd470147757363789, - 64'd30534471519142},
		'{64'd88355216767193600, - 64'd7210717608321972, - 64'd652814047329850, - 64'd74474048717025, 64'd91858913475248672, - 64'd6806001903237092, - 64'd622973704183345, - 64'd72155440125182, 64'd95163132456448672, - 64'd6412774464623528, - 64'd593900038914348, - 64'd69880647819613, 64'd98273569487507344, - 64'd6030841880384146, - 64'd565582022235033, - 64'd67649448246895, 64'd101195823672693504, - 64'd5660010893658376, - 64'd538008559703970, - 64'd65461597775446, 64'd103935397552176256, - 64'd5300088524883438, - 64'd511168501662055, - 64'd63316833651065, 64'd106497697270143200, - 64'd4950882188845119, - 64'd485050652812178, - 64'd61214874927375, 64'd108888032800216368, - 64'd4612199806838576, - 64'd459643781450378, - 64'd59155423371540, 64'd111111618225751072, - 64'd4283849914058110, - 64'd434936628356130, - 64'd57138164345637, 64'd113173572072661216, - 64'd3965641762333352, - 64'd410917915349351, - 64'd55162767664057, 64'd115078917692473632, - 64'd3657385418327684, - 64'd387576353521621, - 64'd53228888427322, 64'd116832583693370816, - 64'd3358891857313212, - 64'd364900651149051, - 64'd51336167832687, 64'd118439404417039040, - 64'd3069973052634992, - 64'd342879521294128, - 64'd49484233961915, 64'd119904120459193856, - 64'd2790442060975596, - 64'd321501689103792, - 64'd47672702546602, 64'd121231379231710912, - 64'd2520113103529546, - 64'd300755898810927, - 64'd45901177711433, 64'd122425735564343952, - 64'd2258801643195464, - 64'd280630920446329, - 64'd44169252695746, 64'd123491652344065504, - 64'd2006324457892246, - 64'd261115556268174, - 64'd42476510553788, 64'd124433501190118432, - 64'd1762499710103830, - 64'd242198646915861, - 64'd40822524834034, 64'd125255563162918528, - 64'd1527147012755594, - 64'd223869077295067, - 64'd39206860237959, 64'd125962029504999408, - 64'd1300087491523733, - 64'd206115782200739, - 64'd37629073258616, 64'd126557002412241056, - 64'd1081143843677293, - 64'd188927751684637, - 64'd36088712799422, 64'd127044495833673088, - 64'd870140393550984, - 64'd172294036173990, - 64'd34585320773506, 64'd127428436298192192, - 64'd666903144745155, - 64'd156203751347696, - 64'd33118432683989, 64'd127712663766581200, - 64'd471259829147740, - 64'd140646082776425, - 64'd31687578185584, 64'd127900932507263808, - 64'd283039952871314, - 64'd125610290332884, - 64'd30292281627854},
		'{64'd88355216767386768, - 64'd7210717608309690, - 64'd652814047329616, - 64'd74474048717007, 64'd91858913475437136, - 64'd6806001903225109, - 64'd622973704183117, - 64'd72155440125165, 64'd95163132456632496, - 64'd6412774464611841, - 64'd593900038914125, - 64'd69880647819597, 64'd98273569487686592, - 64'd6030841880372750, - 64'd565582022234815, - 64'd67649448246879, 64'd101195823672868208, - 64'd5660010893647267, - 64'd538008559703758, - 64'd65461597775430, 64'd103935397552346496, - 64'd5300088524872613, - 64'd511168501661848, - 64'd63316833651049, 64'd106497697270309040, - 64'd4950882188834574, - 64'd485050652811977, - 64'd61214874927360, 64'd108888032800377888, - 64'd4612199806828306, - 64'd459643781450182, - 64'd59155423371526, 64'd111111618225908304, - 64'd4283849914048112, - 64'd434936628355939, - 64'd57138164345623, 64'd113173572072814240, - 64'd3965641762323622, - 64'd410917915349164, - 64'd55162767664043, 64'd115078917692622528, - 64'd3657385418318216, - 64'd387576353521439, - 64'd53228888427309, 64'd116832583693515648, - 64'd3358891857304003, - 64'd364900651148874, - 64'd51336167832674, 64'd118439404417179840, - 64'd3069973052626038, - 64'd342879521293956, - 64'd49484233961902, 64'd119904120459330720, - 64'd2790442060966894, - 64'd321501689103625, - 64'd47672702546590, 64'd121231379231843888, - 64'd2520113103521090, - 64'd300755898810764, - 64'd45901177711421, 64'd122425735564473120, - 64'd2258801643187250, - 64'd280630920446172, - 64'd44169252695734, 64'd123491652344190928, - 64'd2006324457884270, - 64'd261115556268021, - 64'd42476510553776, 64'd124433501190240176, - 64'd1762499710096088, - 64'd242198646915712, - 64'd40822524834023, 64'd125255563163036640, - 64'd1527147012748084, - 64'd223869077294923, - 64'd39206860237948, 64'd125962029505113984, - 64'd1300087491516448, - 64'd206115782200599, - 64'd37629073258605, 64'd126557002412352128, - 64'd1081143843670230, - 64'd188927751684501, - 64'd36088712799412, 64'd127044495833780736, - 64'd870140393544138, - 64'd172294036173858, - 64'd34585320773496, 64'd127428436298296480, - 64'd666903144738522, - 64'd156203751347568, - 64'd33118432683980, 64'd127712663766682176, - 64'd471259829141318, - 64'd140646082776301, - 64'd31687578185574, 64'd127900932507361568, - 64'd283039952865098, - 64'd125610290332764, - 64'd30292281627845}};
	localparam logic signed[63:0] Fbi[0:3][0:99] = '{
		'{- 64'd107703265549738064, - 64'd8947071520977922, 64'd232934047530405, 64'd41073311006417, - 64'd103176552463027872, - 64'd9156640347428454, 64'd203864747109806, 64'd40467587652981, - 64'd98549769089416768, - 64'd9347347755640880, 64'd174926291869582, 64'd39803517402087, - 64'd93832350891096016, - 64'd9519180117281880, 64'd146165341452405, 64'd39083172608701, - 64'd89033732109869584, - 64'd9672155853539060, 64'd117627494402776, 64'd38308686683285, - 64'd84163329879103072, - 64'd9806324880801568, 64'd89357228603024, 64'd37482249497631, - 64'd79230528623918016, - 64'd9921768012283748, 64'd61397844571438, 64'd36606102770485, - 64'd74244664771229408, - 64'd10018596317320144, 64'd33791411671403, 64'd35682535441095, - 64'd69215011790349648, - 64'd10096950440103238, 64'd6578717274732, 64'd34713879038661, - 64'd64150765583986400, - 64'd10156999879674868, - 64'd20200781083337, 64'd33702503055577, - 64'd59061030248547488, - 64'd10198942233017976, - 64'd46509000525631, 64'd32650810332197, - 64'd53954804221733768, - 64'd10223002403127416, - 64'd72309274604807, 64'd31561232460715, - 64'd48840966834455424, - 64'd10229431773966964, - 64'd97566392004763, 64'd30436225215614, - 64'd43728265283145904, - 64'd10218507354244318, - 64'd122246632156539, 64'd29278264017934, - 64'd38625302037577456, - 64'd10190530891956972, - 64'd146317797759052, 64'd28089839440465, - 64'd33540522698301016, - 64'd10145827961679208, - 64'd169749244200350, 64'd26873452760785, - 64'd28482204316844112, - 64'd10084747026574258, - 64'd192511905880381, 64'd25631611568843, - 64'd23458444190805936, - 64'd10007658477125936, - 64'd214578319441481, 64'd24366825435609, - 64'd18477149144990256, - 64'd9914953648590698, - 64'd235922643917893, 64'd23081601649110, - 64'd13546025308714328, - 64'd9807043819174324, - 64'd256520677820646, 64'd21778441023919, - 64'd8672568398431088, - 64'd9684359190937200, - 64'd276349873179018, 64'd20459833789988, - 64'd3864054513799336, - 64'd9547347855428568, - 64'd295389346564595, 64'd19128255566438, 64'd872468545660632, - 64'd9396474746043208, - 64'd313619887128605, 64'd17786163425729, 64'd5530189437183984, - 64'd9232220579083878, - 64'd331023961687728, 64'd16435992053359, 64'd10102540899496720, - 64'd9055080785499432, - 64'd347585716898006, 64'd15080150008005},
		'{64'd107703265549686464, 64'd8947071520974648, - 64'd232934047530462, - 64'd41073311006421, 64'd103176552462974192, 64'd9156640347425048, - 64'd203864747109865, - 64'd40467587652985, 64'd98549769089361104, 64'd9347347755637348, - 64'd174926291869644, - 64'd39803517402091, 64'd93832350891038528, 64'd9519180117278230, - 64'd146165341452470, - 64'd39083172608705, 64'd89033732109810368, 64'd9672155853535304, - 64'd117627494402843, - 64'd38308686683290, 64'd84163329879042272, 64'd9806324880797710, - 64'd89357228603093, - 64'd37482249497635, 64'd79230528623855760, 64'd9921768012279798, - 64'd61397844571508, - 64'd36606102770490, 64'd74244664771165840, 64'd10018596317316110, - 64'd33791411671475, - 64'd35682535441100, 64'd69215011790284872, 64'd10096950440099126, - 64'd6578717274805, - 64'd34713879038666, 64'd64150765583920560, 64'd10156999879670690, 64'd20200781083262, - 64'd33702503055583, 64'd59061030248480696, 64'd10198942233013736, 64'd46509000525554, - 64'd32650810332202, 64'd53954804221666176, 64'd10223002403123124, 64'd72309274604729, - 64'd31561232460721, 64'd48840966834387152, 64'd10229431773962628, 64'd97566392004684, - 64'd30436225215620, 64'd43728265283077064, 64'd10218507354239948, 64'd122246632156459, - 64'd29278264017939, 64'd38625302037508176, 64'd10190530891952574, 64'd146317797758972, - 64'd28089839440471, 64'd33540522698231432, 64'd10145827961674790, 64'd169749244200269, - 64'd26873452760791, 64'd28482204316774328, 64'd10084747026569828, 64'd192511905880300, - 64'd25631611568849, 64'd23458444190736088, 64'd10007658477121504, 64'd214578319441399, - 64'd24366825435615, 64'd18477149144920448, 64'd9914953648586268, 64'd235922643917811, - 64'd23081601649116, 64'd13546025308644696, 64'd9807043819169904, 64'd256520677820564, - 64'd21778441023925, 64'd8672568398361736, 64'd9684359190932798, 64'd276349873178936, - 64'd20459833789994, 64'd3864054513730376, 64'd9547347855424192, 64'd295389346564514, - 64'd19128255566444, - 64'd872468545729080, 64'd9396474746038864, 64'd313619887128524, - 64'd17786163425735, - 64'd5530189437251816, 64'd9232220579079572, 64'd331023961687648, - 64'd16435992053364, - 64'd10102540899563848, 64'd9055080785495172, 64'd347585716897926, - 64'd15080150008011},
		'{- 64'd327914229854852992, - 64'd16132963874025046, - 64'd1038246167410144, - 64'd51020251934053, - 64'd319899697871776704, - 64'd15924753197771214, - 64'd1027886004934731, - 64'd51193749141451, - 64'd311989863798591104, - 64'd15714211612504252, - 64'd1017253638204449, - 64'd51326425925515, - 64'd304185834803758720, - 64'd15501570951755914, - 64'd1006366883742788, - 64'd51419808379449, - 64'd296488604089275968, - 64'd15287055274431814, - 64'd995243022330351, - 64'd51475388318663, - 64'd288899054738239104, - 64'd15070881023600346, - 64'd983898808725565, - 64'd51494623646558, - 64'd281417963483320224, - 64'd14853257184054888, - 64'd972350481349960, - 64'd51478938728343, - 64'd274046004396780480, - 64'd14634385438593302, - 64'd960613771932999, - 64'd51429724772316, - 64'd266783752502675136, - 64'd14414460322961760, - 64'd948703915111656, - 64'd51348340218067, - 64'd259631687311931712, - 64'd14193669379412916, - 64'd936635657980159, - 64'd51236111131066, - 64'd252590196281004288, - 64'd13972193308831394, - 64'd924423269585548, - 64'd51094331603127, - 64'd245659578194833664, - 64'd13750206121382268, - 64'd912080550364871, - 64'd50924264158244, - 64'd238840046474860192, - 64'd13527875285641054, - 64'd899620841520088, - 64'd50727140163322, - 64'd232131732412860224, - 64'd13305361876166310, - 64'd887057034326906, - 64'd50504160243335, - 64'd225534688331392544, - 64'd13082820719478520, - 64'd874401579373997, - 64'd50256494700464, - 64'd219048890671661408, - 64'd12860400538411460, - 64'd861666495729220, - 64'd49985283936770, - 64'd212674243009616960, - 64'd12638244094804652, - 64'd848863380029643, - 64'd49691638879994, - 64'd206410579001130624, - 64'd12416488330507796, - 64'd836003415492366, - 64'd49376641412073, - 64'd200257665257095456, - 64'd12195264506670468, - 64'd823097380843278, - 64'd49041344799975, - 64'd194215204149316032, - 64'd11974698341292420, - 64'd810155659161094, - 64'd48686774128483, - 64'd188282836548062176, - 64'd11754910145012030, - 64'd797188246634127, - 64'd48313926734564, - 64'd182460144492173664, - 64'd11536014955112534, - 64'd784204761227466, - 64'd47923772642960, - 64'd176746653792611072, - 64'd11318122667727552, - 64'd771214451258330, - 64'd47517255002685, - 64'd171141836570357568, - 64'd11101338168229462, - 64'd758226203877556, - 64'd47095290524082, - 64'd165645113729583616, - 64'd10885761459785948, - 64'd745248553455290, - 64'd46658769916138},
		'{64'd327914229854801664, 64'd16132963874021790, 64'd1038246167410088, 64'd51020251934049, 64'd319899697871723264, 64'd15924753197767824, 64'd1027886004934672, 64'd51193749141447, 64'd311989863798535680, 64'd15714211612500738, 64'd1017253638204388, 64'd51326425925511, 64'd304185834803701504, 64'd15501570951752284, 64'd1006366883742724, 64'd51419808379444, 64'd296488604089217024, 64'd15287055274428074, 64'd995243022330285, 64'd51475388318658, 64'd288899054738178496, 64'd15070881023596500, 64'd983898808725497, 64'd51494623646554, 64'd281417963483258144, 64'd14853257184050946, 64'd972350481349890, 64'd51478938728339, 64'd274046004396716960, 64'd14634385438589270, 64'd960613771932928, 64'd51429724772311, 64'd266783752502610304, 64'd14414460322957642, 64'd948703915111582, 64'd51348340218062, 64'd259631687311865600, 64'd14193669379408722, 64'd936635657980084, 64'd51236111131060, 64'd252590196280937088, 64'd13972193308827128, 64'd924423269585471, 64'd51094331603121, 64'd245659578194765408, 64'd13750206121377934, 64'd912080550364793, 64'd50924264158238, 64'd238840046474790976, 64'd13527875285636658, 64'd899620841520008, 64'd50727140163316, 64'd232131732412790144, 64'd13305361876161860, 64'd887057034326825, 64'd50504160243330, 64'd225534688331321664, 64'd13082820719474018, 64'd874401579373915, 64'd50256494700458, 64'd219048890671589760, 64'd12860400538406916, 64'd861666495729137, 64'd49985283936764, 64'd212674243009544736, 64'd12638244094800064, 64'd848863380029560, 64'd49691638879988, 64'd206410579001057824, 64'd12416488330503172, 64'd836003415492282, 64'd49376641412067, 64'd200257665257022144, 64'd12195264506665812, 64'd823097380843194, 64'd49041344799968, 64'd194215204149242304, 64'd11974698341287738, 64'd810155659161008, 64'd48686774128477, 64'd188282836547988064, 64'd11754910145007324, 64'd797188246634041, 64'd48313926734557, 64'd182460144492099264, 64'd11536014955107808, 64'd784204761227379, 64'd47923772642954, 64'd176746653792536448, 64'd11318122667722810, 64'd771214451258244, 64'd47517255002679, 64'd171141836570282784, 64'd11101338168224710, 64'd758226203877469, 64'd47095290524076, 64'd165645113729508704, 64'd10885761459781186, 64'd745248553455202, 64'd46658769916132}};
	localparam logic signed[63:0] hf[0:1199] = {64'd3920895148032, - 64'd2763445504, - 64'd3587446528, 64'd4984890, 64'd3918132150272, - 64'd8286441984, - 64'd3577147648, 64'd14935367, 64'd3912610611200, - 64'd13797770240, - 64'd3556578816, 64'd24828730, 64'd3904337608704, - 64'd19289686016, - 64'd3525795840, 64'd34628620, 64'd3893325463552, - 64'd24754487296, - 64'd3484879104, 64'd44300172, 64'd3879589117952, - 64'd30184531968, - 64'd3433933312, 64'd53810032, 64'd3863147970560, - 64'd35572252672, - 64'd3373086976, 64'd63126368, 64'd3844025090048, - 64'd40910168064, - 64'd3302491136, 64'd72218896, 64'd3822247215104, - 64'd46190915584, - 64'd3222318592, 64'd81058880, 64'd3797844754432, - 64'd51407228928, - 64'd3132763136, 64'd89619136, 64'd3770851786752, - 64'd56551993344, - 64'd3034038528, 64'd97874048, 64'd3741305798656, - 64'd61618237440, - 64'd2926377728, 64'd105799568, 64'd3709247946752, - 64'd66599137280, - 64'd2810031616, 64'd113373200, 64'd3674722009088, - 64'd71488045056, - 64'd2685268736, 64'd120574040, 64'd3637776220160, - 64'd76278505472, - 64'd2552373504, 64'd127382712, 64'd3598460911616, - 64'd80964231168, - 64'd2411645696, 64'd133781400, 64'd3556830347264, - 64'd85539176448, - 64'd2263399424, 64'd139753840, 64'd3512941412352, - 64'd89997467648, - 64'd2107962496, 64'd145285280, 64'd3466853351424, - 64'd94333476864, - 64'd1945674752, 64'd150362496, 64'd3418629079040, - 64'd98541805568, - 64'd1776887552, 64'd154973776, 64'd3368333606912, - 64'd102617292800, - 64'd1601962880, 64'd159108848, 64'd3316034830336, - 64'd106555015168, - 64'd1421272064, 64'd162758960, 64'd3261802479616, - 64'd110350319616, - 64'd1235195008, 64'd165916736, 64'd3205708906496, - 64'd113998798848, - 64'd1044119040, 64'd168576256, 64'd3147828822016, - 64'd117496307712, - 64'd848438400, 64'd170732992, 64'd3088238247936, - 64'd120838995968, - 64'd648552768, 64'd172383744, 64'd3027016089600, - 64'd124023259136, - 64'd444866688, 64'd173526688, 64'd2964242038784, - 64'd127045787648, - 64'd237788400, 64'd174161264, 64'd2899997884416, - 64'd129903550464, - 64'd27729112, 64'd174288224, 64'd2834366464000, - 64'd132593795072, 64'd184897952, 64'd173909488, 64'd2767432187904, - 64'd135114063872, 64'd399678464, 64'd173028256, 64'd2699281039360, - 64'd137462185984, 64'd616197888, 64'd171648848, 64'd2629999001600, - 64'd139636293632, 64'd834042176, 64'd169776720, 64'd2559673892864, - 64'd141634748416, 64'd1052798720, 64'd167418416, 64'd2488393793536, - 64'd143456288768, 64'd1272057344, 64'd164581536, 64'd2416247308288, - 64'd145099898880, 64'd1491410560, 64'd161274688, 64'd2343323828224, - 64'd146564808704, 64'd1710454912, 64'd157507440, 64'd2269712482304, - 64'd147850625024, 64'd1928791424, 64'd153290288, 64'd2195503054848, - 64'd148957151232, 64'd2146026496, 64'd148634624, 64'd2120785068032, - 64'd149884534784, 64'd2361772032, 64'd143552672, 64'd2045648306176, - 64'd150633152512, 64'd2575647488, 64'd138057456, 64'd1970181636096, - 64'd151203692544, 64'd2787278336, 64'd132162728, 64'd1894474055680, - 64'd151597088768, 64'd2996299264, 64'd125882992, 64'd1818613907456, - 64'd151814569984, 64'd3202352384, 64'd119233376, 64'd1742688616448, - 64'd151857577984, 64'd3405089792, 64'd112229640, 64'd1666785083392, - 64'd151727833088, 64'd3604172288, 64'd104888120, 64'd1590989160448, - 64'd151427334144, 64'd3799271680, 64'd97225680, 64'd1515385782272, - 64'd150958276608, 64'd3990069760, 64'd89259656, 64'd1440058572800, - 64'd150323101696, 64'd4176259584, 64'd81007824, 64'd1365089976320, - 64'd149524512768, 64'd4357545984, 64'd72488360, 64'd1290560864256, - 64'd148565409792, 64'd4533644800, 64'd63719772, 64'd1216550797312, - 64'd147448905728, 64'd4704285696, 64'd54720884, 64'd1143137632256, - 64'd146178310144, 64'd4869209600, 64'd45510776, 64'd1070397587456, - 64'd144757178368, 64'd5028170752, 64'd36108744, 64'd998404980736, - 64'd143189213184, 64'd5180936704, 64'd26534250, 64'd927232229376, - 64'd141478297600, 64'd5327288320, 64'd16806892, 64'd856949784576, - 64'd139628527616, 64'd5467019776, 64'd6946355, 64'd787626131456, - 64'd137644146688, 64'd5599940608, - 64'd3027632, 64'd719327330304, - 64'd135529529344, 64'd5725872640, - 64'd13095330, 64'd652117540864, - 64'd133289222144, 64'd5844652032, - 64'd23237034, 64'd586058301440, - 64'd130927910912, 64'd5956130816, - 64'd33433110, 64'd521208987648, - 64'd128450404352, 64'd6060173824, - 64'd43664036, 64'd457626451968, - 64'd125861625856, 64'd6156660736, - 64'd53910432, 64'd395365056512, - 64'd123166621696, 64'd6245485568, - 64'd64153100, 64'd334476673024, - 64'd120370511872, 64'd6326557184, - 64'd74373064, 64'd275010551808, - 64'd117478539264, 64'd6399797760, - 64'd84551600, 64'd217013239808, - 64'd114496012288, 64'd6465145856, - 64'd94670248, 64'd160528728064, - 64'd111428296704, 64'd6522552320, - 64'd104710888, 64'd105598238720, - 64'd108280840192, 64'd6571982848, - 64'd114655736, 64'd52260270080, - 64'd105059131392, 64'd6613417472, - 64'd124487368, 64'd550564480, - 64'd101768708096, 64'd6646850048, - 64'd134188784, - 64'd49497907200, - 64'd98415132672, 64'd6672287232, - 64'd143743392, - 64'd97854971904, - 64'd95003992064, 64'd6689750528, - 64'd153135072, - 64'd144493232128, - 64'd91540897792, 64'd6699274240, - 64'd162348160, - 64'd189388128256, - 64'd88031444992, 64'd6700904960, - 64'd171367520, - 64'd232517894144, - 64'd84481245184, 64'd6694703104, - 64'd180178512, - 64'd273863507968, - 64'd80895877120, 64'd6680741376, - 64'd188767040, - 64'd313408815104, - 64'd77280911360, 64'd6659104768, - 64'd197119584, - 64'd351140413440, - 64'd73641885696, 64'd6629889024, - 64'd205223200, - 64'd387047620608, - 64'd69984296960, 64'd6593203200, - 64'd213065504, - 64'd421122506752, - 64'd66313576448, 64'd6549166592, - 64'd220634768, - 64'd453359894528, - 64'd62635130880, 64'd6497910272, - 64'd227919840, - 64'd483757228032, - 64'd58954276864, 64'd6439574016, - 64'd234910240, - 64'd512314638336, - 64'd55276269568, 64'd6374309376, - 64'd241596096, - 64'd539034845184, - 64'd51606282240, 64'd6302277632, - 64'd247968224, - 64'd563923124224, - 64'd47949410304, 64'd6223648256, - 64'd254018064, - 64'd586987274240, - 64'd44310642688, 64'd6138600448, - 64'd259737728, - 64'd608237584384, - 64'd40694874112, 64'd6047321600, - 64'd265120032, - 64'd627686768640, - 64'd37106892800, 64'd5950007296, - 64'd270158432, - 64'd645349900288, - 64'd33551376384, 64'd5846860800, - 64'd274847072, - 64'd661244346368, - 64'd30032877568, 64'd5738092032, - 64'd279180768, - 64'd675389702144, - 64'd26555826176, 64'd5623918592, - 64'd283155040, - 64'd687807791104, - 64'd23124529152, 64'd5504562688, - 64'd286766048, - 64'd698522533888, - 64'd19743150080, 64'd5380253696, - 64'd290010656, - 64'd707559882752, - 64'd16415717376, 64'd5251225600, - 64'd292886368, - 64'd714947887104, - 64'd13146114048, 64'd5117718016, - 64'd295391392, - 64'd720716300288, - 64'd9938075648, 64'd4979973632, - 64'd297524544, - 64'd724896776192, - 64'd6795185152, 64'd4838239744, - 64'd299285376, - 64'd727522869248, - 64'd3720871424, 64'd4692767232, - 64'd300673984, - 64'd728629641216, - 64'd718402880, 64'd4543809536, - 64'd301691168, - 64'd728253792256, 64'd2209112576, 64'd4391622656, - 64'd302338336, - 64'd726433529856, 64'd5058731520, 64'd4236464640, - 64'd302617536, - 64'd723208503296, 64'd7827677696, 64'd4078595328, - 64'd302531328, - 64'd718619738112, 64'd10513341440, 64'd3918274816, - 64'd302082976, - 64'd712709439488, 64'd13113285632, 64'd3755764480, - 64'd301276256, - 64'd705521123328, 64'd15625242624, 64'd3591326208, - 64'd300115520, - 64'd697099223040, 64'd18047119360, 64'd3425220608, - 64'd298605664, - 64'd687489286144, 64'd20376993792, 64'd3257708288, - 64'd296752064, - 64'd676737843200, 64'd22613118976, 64'd3089048576, - 64'd294560736, - 64'd664892080128, 64'd24753920000, 64'd2919499520, - 64'd292038048, - 64'd652000034816, 64'd26798000128, 64'd2749316608, - 64'd289190944, - 64'd638110400512, 64'd28744130560, 64'd2578753536, - 64'd286026784, - 64'd623272394752, 64'd30591258624, 64'd2408060928, - 64'd282553408, - 64'd607535759360, 64'd32338505728, 64'd2237486336, - 64'd278778976, - 64'd590950694912, 64'd33985155072, 64'd2067274112, - 64'd274712192, - 64'd573567467520, 64'd35530665984, 64'd1897664256, - 64'd270361984, - 64'd555436933120, 64'd36974665728, 64'd1728892928, - 64'd265737808, - 64'd536609783808, 64'd38316945408, 64'd1561191680, - 64'd260849328, - 64'd517136941056, 64'd39557451776, 64'd1394787200, - 64'd255706560, - 64'd497069260800, 64'd40696303616, 64'd1229901184, - 64'd250319824, - 64'd476457533440, 64'd41733771264, 64'd1066749632, - 64'd244699744, - 64'd455352320000, 64'd42670284800, 64'd905542912, - 64'd238857120, - 64'd433803984896, 64'd43506413568, 64'd746485440, - 64'd232803056, - 64'd411862532096, 64'd44242890752, 64'd589775296, - 64'd226548832, - 64'd389577572352, 64'd44880584704, 64'd435604288, - 64'd220105888, - 64'd366998224896, 64'd45420507136, 64'd284157280, - 64'd213485872, - 64'd344173150208, 64'd45863813120, 64'd135612352, - 64'd206700560, - 64'd321150320640, 64'd46211780608, - 64'd9859543, - 64'd199761840, - 64'd297977020416, 64'd46465826816, - 64'd152094736, - 64'd192681680, - 64'd274699894784, 64'd46627483648, - 64'd290937024, - 64'd185472160, - 64'd251364671488, 64'd46698405888, - 64'd426237760, - 64'd178145408, - 64'd228016308224, 64'd46680375296, - 64'd557856064, - 64'd170713552, - 64'd204698812416, 64'd46575267840, - 64'd685658880, - 64'd163188784, - 64'd181455224832, 64'd46385074176, - 64'd809521088, - 64'd155583232, - 64'd158327570432, 64'd46111883264, - 64'd929325632, - 64'd147909040, - 64'd135356817408, 64'd45757886464, - 64'd1044963584, - 64'd140178272, - 64'd112582778880, 64'd45325357056, - 64'd1156334208, - 64'd132402944, - 64'd90044153856, 64'd44816658432, - 64'd1263344768, - 64'd124594992, - 64'd67778412544, 64'd44234235904, - 64'd1365911168, - 64'd116766208, - 64'd45821788160, 64'd43580604416, - 64'd1463957248, - 64'd108928312, - 64'd24209246208, 64'd42858356736, - 64'd1557415168, - 64'd101092824, - 64'd2974428672, 64'd42070142976, - 64'd1646225536, - 64'd93271160, 64'd17850353664, 64'd41218678784, - 64'd1730336896, - 64'd85474520, 64'd38234165248, 64'd40306724864, - 64'd1809705984, - 64'd77713928, 64'd58147467264, 64'd39337099264, - 64'd1884298112, - 64'd70000208, 64'd77562126336, 64'd38312656896, - 64'd1954086144, - 64'd62343932, 64'd96451469312, 64'd37236293632, - 64'd2019051008, - 64'd54755468, 64'd114790252544, 64'd36110934016, - 64'd2079181952, - 64'd47244916, 64'd132554727424, 64'd34939535360, - 64'd2134475520, - 64'd39822112, 64'd149722611712, 64'd33725071360, - 64'd2184935936, - 64'd32496616, 64'd166273122304, 64'd32470532096, - 64'd2230575616, - 64'd25277704, 64'd182186967040, 64'd31178921984, - 64'd2271413760, - 64'd18174346, 64'd197446352896, 64'd29853249536, - 64'd2307476992, - 64'd11195207, 64'd212035026944, 64'd28496527360, - 64'd2338799104, - 64'd4348626, 64'd225938210816, 64'd27111757824, - 64'd2365421056, 64'd2357381, 64'd239142617088, 64'd25701941248, - 64'd2387390208, 64'd8915142, 64'd251636465664, 64'd24270059520, - 64'd2404760576, 64'd15317325, 64'd263409483776, 64'd22819080192, - 64'd2417593088, 64'd21556954, 64'd274452856832, 64'd21351946240, - 64'd2425954048, 64'd27627412, 64'd284759228416, 64'd19871571968, - 64'd2429916672, 64'd33522442, 64'd294322700288, 64'd18380845056, - 64'd2429559296, 64'd39236160, 64'd303138832384, 64'd16882610176, - 64'd2424966144, 64'd44763060, 64'd311204511744, 64'd15379678208, - 64'd2416226560, 64'd50098004, 64'd318518165504, 64'd13874812928, - 64'd2403435264, 64'd55236240, 64'd325079465984, 64'd12370733056, - 64'd2386691840, 64'd60173392, 64'd330889494528, 64'd10870104064, - 64'd2366100224, 64'd64905476, 64'd335950577664, 64'd9375537152, - 64'd2341769216, 64'd69428888, 64'd340266450944, 64'd7889585664, - 64'd2313811200, 64'd73740416, 64'd343842029568, 64'd6414739968, - 64'd2282343168, 64'd77837216, 64'd346683441152, 64'd4953428480, - 64'd2247484928, 64'd81716832, 64'd348798091264, 64'd3508009728, - 64'd2209360640, 64'd85377208, 64'd350194499584, 64'd2080774016, - 64'd2168096512, 64'd88816648, 64'd350882267136, 64'd673937472, - 64'd2123822848, 64'd92033824, 64'd350872174592, - 64'd710358208, - 64'd2076671616, 64'd95027808, 64'd350176018432, - 64'd2070049152, - 64'd2026777600, 64'd97798024, 64'd348806545408, - 64'd3403151104, - 64'd1974277376, 64'd100344256, 64'd346777616384, - 64'd4707761152, - 64'd1919309952, 64'd102666648, 64'd344103845888, - 64'd5982059520, - 64'd1862015232, 64'd104765704, 64'd340800897024, - 64'd7224311808, - 64'd1802534912, 64'd106642272, 64'd336885153792, - 64'd8432869888, - 64'd1741011712, 64'd108297536, 64'd332373884928, - 64'd9606172672, - 64'd1677589120, 64'd109733016, 64'd327285112832, - 64'd10742748160, - 64'd1612411136, 64'd110950552, 64'd321637482496, - 64'd11841213440, - 64'd1545622144, 64'd111952312, 64'd315450458112, - 64'd12900276224, - 64'd1477366784, 64'd112740760, 64'd308743995392, - 64'd13918737408, - 64'd1407789440, 64'd113318664, 64'd301538672640, - 64'd14895484928, - 64'd1337033984, 64'd113689088, 64'd293855625216, - 64'd15829501952, - 64'd1265243904, 64'd113855368, 64'd285716447232, - 64'd16719862784, - 64'd1192561792, 64'd113821120, 64'd277143191552, - 64'd17565732864, - 64'd1119129088, 64'd113590208, 64'd268158255104, - 64'd18366367744, - 64'd1045086016, 64'd113166760, 64'd258784460800, - 64'd19121117184, - 64'd970571456, 64'd112555144, 64'd249044877312, - 64'd19829422080, - 64'd895722432, 64'd111759944, 64'd238962851840, - 64'd20490811392, - 64'd820674112, 64'd110785976, 64'd228561944576, - 64'd21104902144, - 64'd745559744, 64'd109638248, 64'd217865879552, - 64'd21671403520, - 64'd670510080, 64'd108321976, 64'd206898511872, - 64'd22190108672, - 64'd595653696, 64'd106842552, 64'd195683762176, - 64'd22660902912, - 64'd521116320, 64'd105205544, 64'd184245600256, - 64'd23083747328, - 64'd447021088, 64'd103416680, 64'd172607995904, - 64'd23458697216, - 64'd373488128, 64'd101481824, 64'd160794869760, - 64'd23785879552, - 64'd300634528, 64'd99407000, 64'd148830044160, - 64'd24065511424, - 64'd228574128, 64'd97198328, 64'd136737234944, - 64'd24297881600, - 64'd157417440, 64'd94862056, 64'd124539977728, - 64'd24483358720, - 64'd87271464, 64'd92404536, 64'd112261619712, - 64'd24622387200, - 64'd18239634, 64'd89832192, 64'd99925254144, - 64'd24715481088, 64'd49578332, 64'd87151536, 64'd87553695744, - 64'd24763226112, 64'd116086544, 64'd84369136, 64'd75169472512, - 64'd24766281728, 64'd181192992, 64'd81491624, 64'd62794747904, - 64'd24725364736, 64'd244809696, 64'd78525664, 64'd50451308544, - 64'd24641265664, 64'd306852736, 64'd75477936, 64'd38160543744, - 64'd24514826240, 64'd367242272, 64'd72355168, 64'd25943390208, - 64'd24346955776, 64'd425902784, 64'd69164072, 64'd13820332032, - 64'd24138616832, 64'd482762944, 64'd65911356, 64'd1811350400, - 64'd23890825216, 64'd537755776, 64'd62603716, - 64'd10064093184, - 64'd23604645888, 64'd590818496, 64'd59247820, - 64'd21787082752, - 64'd23281199104, 64'd641892992, 64'd55850300, - 64'd33339271168, - 64'd22921641984, 64'd690925248, 64'd52417744, - 64'd44702904320, - 64'd22527182848, 64'd737865792, 64'd48956668, - 64'd55860842496, - 64'd22099064832, 64'd782669696, 64'd45473540, - 64'd66796572672, - 64'd21638572032, 64'd825296256, 64'd41974736, - 64'd77494239232, - 64'd21147019264, 64'd865709248, 64'd38466552, - 64'd87938637824, - 64'd20625756160, 64'd903876928, 64'd34955184, - 64'd98115272704, - 64'd20076163072, 64'd939771840, 64'd31446734, - 64'd108010307584, - 64'd19499638784, 64'd973370944, 64'd27947182, - 64'd117610659840, - 64'd18897614848, 64'd1004655424, 64'd24462388, - 64'd126903918592, - 64'd18271537152, 64'd1033610880, 64'd20998092, - 64'd135878426624, - 64'd17622872064, 64'd1060227008, 64'd17559890, - 64'd144523264000, - 64'd16953097216, 64'd1084497792, 64'd14153241, - 64'd152828248064, - 64'd16263705600, 64'd1106421120, 64'd10783452, - 64'd160783958016, - 64'd15556200448, 64'd1125999232, 64'd7455676, - 64'd168381677568, - 64'd14832087040, 64'd1143238144, 64'd4174906, - 64'd175613526016, - 64'd14092879872, 64'd1158147712, 64'd945966, - 64'd182472294400, - 64'd13340089344, 64'd1170741760, - 64'd2226493, - 64'd188951592960, - 64'd12575229952, 64'd1181037824, - 64'd5337993, - 64'd195045769216, - 64'd11799806976, 64'd1189057024, - 64'd8384241, - 64'd200749891584, - 64'd11015324672, 64'd1194823808, - 64'd11361127, - 64'd206059831296, - 64'd10223272960, 64'd1198366464, - 64'd14264733, - 64'd210972147712, - 64'd9425134592, 64'd1199716352, - 64'd17091330, - 64'd215484186624, - 64'd8622377984, 64'd1198908160, - 64'd19837388, - 64'd219593998336, - 64'd7816452608, 64'd1195979520, - 64'd22499570, - 64'd223300354048, - 64'd7008794112, 64'd1190971136, - 64'd25074746, - 64'd226602745856, - 64'd6200815104, 64'd1183926656, - 64'd27559984, - 64'd229501353984, - 64'd5393906688, 64'd1174892416, - 64'd29952556, - 64'd231997046784, - 64'd4589435904, 64'd1163917312, - 64'd32249940, - 64'd234091413504, - 64'd3788742912, 64'd1151052928, - 64'd34449816, - 64'd235786649600, - 64'd2993140224, 64'd1136353024, - 64'd36550072, - 64'd237085605888, - 64'd2203910400, 64'd1119873664, - 64'd38548808, - 64'd237991821312, - 64'd1422304256, 64'd1101672960, - 64'd40444320, - 64'd238509391872, - 64'd649539328, 64'd1081811200, - 64'd42235112, - 64'd238643036160, 64'd113201360, 64'd1060350080, - 64'd43919896, - 64'd238398046208, 64'd864771136, 64'd1037353472, - 64'd45497580, - 64'd237780303872, 64'd1604060800, 64'd1012886464, - 64'd46967280, - 64'd236796215296, 64'd2329999872, 64'd987015808, - 64'd48328308, - 64'd235452710912, 64'd3041558016, 64'd959809408, - 64'd49580176, - 64'd233757212672, 64'd3737746176, 64'd931336320, - 64'd50722580, - 64'd231717683200, 64'd4417616896, 64'd901666624, - 64'd51755424, - 64'd229342461952, 64'd5080265728, 64'd870871360, - 64'd52678784, - 64'd226640429056, 64'd5724833280, 64'd839022144, - 64'd53492940, - 64'd223620792320, 64'd6350503424, 64'd806191424, - 64'd54198332, - 64'd220293201920, 64'd6956505600, 64'd772451904, - 64'd54795596, - 64'd216667684864, 64'd7542115840, 64'd737876800, - 64'd55285532, - 64'd212754595840, 64'd8106655744, 64'd702539392, - 64'd55669116, - 64'd208564633600, 64'd8649493504, 64'd666513216, - 64'd55947480, - 64'd204108808192, 64'd9170045952, 64'd629871616, - 64'd56121928, - 64'd199398391808, 64'd9667774464, 64'd592687872, - 64'd56193908, - 64'd194444918784, 64'd10142189568, 64'd555034944, - 64'd56165024, - 64'd189260169216, 64'd10592849920, 64'd516985344, - 64'd56037028, - 64'd183856103424, 64'd11019360256, 64'd478611136, - 64'd55811808, - 64'd178244894720, 64'd11421373440, 64'd439983712, - 64'd55491384, - 64'd172438863872, 64'd11798588416, 64'd401173696, - 64'd55077908, - 64'd166450479104, 64'd12150753280, 64'd362250944, - 64'd54573656, - 64'd160292323328, 64'd12477660160, 64'd323284256, - 64'd53981016, - 64'd153977044992, 64'd12779149312, 64'd284341408, - 64'd53302488, - 64'd147517423616, 64'd13055105024, 64'd245489072, - 64'd52540680, - 64'd140926222336, 64'd13305457664, 64'd206792592, - 64'd51698296, - 64'd134216237056, 64'd13530182656, 64'd168316000, - 64'd50778136, - 64'd127400304640, 64'd13729299456, 64'd130121920, - 64'd49783076, - 64'd120491196416, 64'd13902867456, 64'd92271440, - 64'd48716084, - 64'd113501675520, 64'd14050993152, 64'd54824076, - 64'd47580192, - 64'd106444423168, 64'd14173821952, 64'd17837676, - 64'd46378508, - 64'd99332038656, 64'd14271538176, - 64'd18631644, - 64'd45114188, - 64'd92177031168, 64'd14344369152, - 64'd54529576, - 64'd43790452, - 64'd84991770624, 64'd14392578048, - 64'd89803664, - 64'd42410568, - 64'd77788504064, 64'd14416467968, - 64'd124403384, - 64'd40977836, - 64'd70579306496, 64'd14416375808, - 64'd158280192, - 64'd39495604, - 64'd63376064512, 64'd14392675328, - 64'd191387552, - 64'd37967240, - 64'd56190496768, 64'd14345773056, - 64'd223681008, - 64'd36396140, - 64'd49034088448, 64'd14276109312, - 64'd255118208, - 64'd34785712, - 64'd41918103552, 64'd14184155136, - 64'd285658976, - 64'd33139376, - 64'd34853564416, 64'd14070413312, - 64'd315265312, - 64'd31460558, - 64'd27851235328, 64'd13935413248, - 64'd343901376, - 64'd29752682, - 64'd20921602048, 64'd13779713024, - 64'd371533664, - 64'd28019164, - 64'd14074874880, 64'd13603896320, - 64'd398130784, - 64'd26263408, - 64'd7320958464, 64'd13408571392, - 64'd423663776, - 64'd24488800, - 64'd669450048, 64'd13194371072, - 64'd448105888, - 64'd22698702, 64'd5870374912, 64'd12961948672, - 64'd471432608, - 64'd20896444, 64'd12289572864, 64'd12711977984, - 64'd493621792, - 64'd19085330, 64'd18579542016, 64'd12445151232, - 64'd514653600, - 64'd17268614, 64'd24732033024, 64'd12162180096, - 64'd534510400, - 64'd15449513, 64'd30739152896, 64'd11863788544, - 64'd553176960, - 64'd13631193, 64'd36593373184, 64'd11550717952, - 64'd570640256, - 64'd11816766};
	localparam logic signed[63:0] hb[0:1199] = {64'd3920895148032, 64'd2763445504, - 64'd3587446528, - 64'd4984890, 64'd3918132150272, 64'd8286441984, - 64'd3577147648, - 64'd14935367, 64'd3912610611200, 64'd13797770240, - 64'd3556578816, - 64'd24828730, 64'd3904337608704, 64'd19289686016, - 64'd3525795840, - 64'd34628620, 64'd3893325463552, 64'd24754487296, - 64'd3484879104, - 64'd44300172, 64'd3879589117952, 64'd30184531968, - 64'd3433933312, - 64'd53810032, 64'd3863147970560, 64'd35572252672, - 64'd3373086976, - 64'd63126368, 64'd3844025090048, 64'd40910168064, - 64'd3302491136, - 64'd72218896, 64'd3822247215104, 64'd46190915584, - 64'd3222318592, - 64'd81058880, 64'd3797844754432, 64'd51407228928, - 64'd3132763136, - 64'd89619136, 64'd3770851786752, 64'd56551993344, - 64'd3034038528, - 64'd97874048, 64'd3741305798656, 64'd61618237440, - 64'd2926377728, - 64'd105799568, 64'd3709247946752, 64'd66599137280, - 64'd2810031616, - 64'd113373200, 64'd3674722009088, 64'd71488045056, - 64'd2685268736, - 64'd120574040, 64'd3637776220160, 64'd76278505472, - 64'd2552373504, - 64'd127382712, 64'd3598460911616, 64'd80964231168, - 64'd2411645696, - 64'd133781400, 64'd3556830347264, 64'd85539176448, - 64'd2263399424, - 64'd139753840, 64'd3512941412352, 64'd89997467648, - 64'd2107962496, - 64'd145285280, 64'd3466853351424, 64'd94333476864, - 64'd1945674752, - 64'd150362496, 64'd3418629079040, 64'd98541805568, - 64'd1776887552, - 64'd154973776, 64'd3368333606912, 64'd102617292800, - 64'd1601962880, - 64'd159108848, 64'd3316034830336, 64'd106555015168, - 64'd1421272064, - 64'd162758960, 64'd3261802479616, 64'd110350319616, - 64'd1235195008, - 64'd165916736, 64'd3205708906496, 64'd113998798848, - 64'd1044119040, - 64'd168576256, 64'd3147828822016, 64'd117496307712, - 64'd848438400, - 64'd170732992, 64'd3088238247936, 64'd120838995968, - 64'd648552768, - 64'd172383744, 64'd3027016089600, 64'd124023259136, - 64'd444866688, - 64'd173526688, 64'd2964242038784, 64'd127045787648, - 64'd237788400, - 64'd174161264, 64'd2899997884416, 64'd129903550464, - 64'd27729112, - 64'd174288224, 64'd2834366464000, 64'd132593795072, 64'd184897952, - 64'd173909488, 64'd2767432187904, 64'd135114063872, 64'd399678464, - 64'd173028256, 64'd2699281039360, 64'd137462185984, 64'd616197888, - 64'd171648848, 64'd2629999001600, 64'd139636293632, 64'd834042176, - 64'd169776720, 64'd2559673892864, 64'd141634748416, 64'd1052798720, - 64'd167418416, 64'd2488393793536, 64'd143456288768, 64'd1272057344, - 64'd164581536, 64'd2416247308288, 64'd145099898880, 64'd1491410560, - 64'd161274688, 64'd2343323828224, 64'd146564808704, 64'd1710454912, - 64'd157507440, 64'd2269712482304, 64'd147850625024, 64'd1928791424, - 64'd153290288, 64'd2195503054848, 64'd148957151232, 64'd2146026496, - 64'd148634624, 64'd2120785068032, 64'd149884534784, 64'd2361772032, - 64'd143552672, 64'd2045648306176, 64'd150633152512, 64'd2575647488, - 64'd138057456, 64'd1970181636096, 64'd151203692544, 64'd2787278336, - 64'd132162728, 64'd1894474055680, 64'd151597088768, 64'd2996299264, - 64'd125882992, 64'd1818613907456, 64'd151814569984, 64'd3202352384, - 64'd119233376, 64'd1742688616448, 64'd151857577984, 64'd3405089792, - 64'd112229640, 64'd1666785083392, 64'd151727833088, 64'd3604172288, - 64'd104888120, 64'd1590989160448, 64'd151427334144, 64'd3799271680, - 64'd97225680, 64'd1515385782272, 64'd150958276608, 64'd3990069760, - 64'd89259656, 64'd1440058572800, 64'd150323101696, 64'd4176259584, - 64'd81007824, 64'd1365089976320, 64'd149524512768, 64'd4357545984, - 64'd72488360, 64'd1290560864256, 64'd148565409792, 64'd4533644800, - 64'd63719772, 64'd1216550797312, 64'd147448905728, 64'd4704285696, - 64'd54720884, 64'd1143137632256, 64'd146178310144, 64'd4869209600, - 64'd45510776, 64'd1070397587456, 64'd144757178368, 64'd5028170752, - 64'd36108744, 64'd998404980736, 64'd143189213184, 64'd5180936704, - 64'd26534250, 64'd927232229376, 64'd141478297600, 64'd5327288320, - 64'd16806892, 64'd856949784576, 64'd139628527616, 64'd5467019776, - 64'd6946355, 64'd787626131456, 64'd137644146688, 64'd5599940608, 64'd3027632, 64'd719327330304, 64'd135529529344, 64'd5725872640, 64'd13095330, 64'd652117540864, 64'd133289222144, 64'd5844652032, 64'd23237034, 64'd586058301440, 64'd130927910912, 64'd5956130816, 64'd33433110, 64'd521208987648, 64'd128450404352, 64'd6060173824, 64'd43664036, 64'd457626451968, 64'd125861625856, 64'd6156660736, 64'd53910432, 64'd395365056512, 64'd123166621696, 64'd6245485568, 64'd64153100, 64'd334476673024, 64'd120370511872, 64'd6326557184, 64'd74373064, 64'd275010551808, 64'd117478539264, 64'd6399797760, 64'd84551600, 64'd217013239808, 64'd114496012288, 64'd6465145856, 64'd94670248, 64'd160528728064, 64'd111428296704, 64'd6522552320, 64'd104710888, 64'd105598238720, 64'd108280840192, 64'd6571982848, 64'd114655736, 64'd52260270080, 64'd105059131392, 64'd6613417472, 64'd124487368, 64'd550564480, 64'd101768708096, 64'd6646850048, 64'd134188784, - 64'd49497907200, 64'd98415132672, 64'd6672287232, 64'd143743392, - 64'd97854971904, 64'd95003992064, 64'd6689750528, 64'd153135072, - 64'd144493232128, 64'd91540897792, 64'd6699274240, 64'd162348160, - 64'd189388128256, 64'd88031444992, 64'd6700904960, 64'd171367520, - 64'd232517894144, 64'd84481245184, 64'd6694703104, 64'd180178512, - 64'd273863507968, 64'd80895877120, 64'd6680741376, 64'd188767040, - 64'd313408815104, 64'd77280911360, 64'd6659104768, 64'd197119584, - 64'd351140413440, 64'd73641885696, 64'd6629889024, 64'd205223200, - 64'd387047620608, 64'd69984296960, 64'd6593203200, 64'd213065504, - 64'd421122506752, 64'd66313576448, 64'd6549166592, 64'd220634768, - 64'd453359894528, 64'd62635130880, 64'd6497910272, 64'd227919840, - 64'd483757228032, 64'd58954276864, 64'd6439574016, 64'd234910240, - 64'd512314638336, 64'd55276269568, 64'd6374309376, 64'd241596096, - 64'd539034845184, 64'd51606282240, 64'd6302277632, 64'd247968224, - 64'd563923124224, 64'd47949410304, 64'd6223648256, 64'd254018064, - 64'd586987274240, 64'd44310642688, 64'd6138600448, 64'd259737728, - 64'd608237584384, 64'd40694874112, 64'd6047321600, 64'd265120032, - 64'd627686768640, 64'd37106892800, 64'd5950007296, 64'd270158432, - 64'd645349900288, 64'd33551376384, 64'd5846860800, 64'd274847072, - 64'd661244346368, 64'd30032877568, 64'd5738092032, 64'd279180768, - 64'd675389702144, 64'd26555826176, 64'd5623918592, 64'd283155040, - 64'd687807791104, 64'd23124529152, 64'd5504562688, 64'd286766048, - 64'd698522533888, 64'd19743150080, 64'd5380253696, 64'd290010656, - 64'd707559882752, 64'd16415717376, 64'd5251225600, 64'd292886368, - 64'd714947887104, 64'd13146114048, 64'd5117718016, 64'd295391392, - 64'd720716300288, 64'd9938075648, 64'd4979973632, 64'd297524544, - 64'd724896776192, 64'd6795185152, 64'd4838239744, 64'd299285376, - 64'd727522869248, 64'd3720871424, 64'd4692767232, 64'd300673984, - 64'd728629641216, 64'd718402880, 64'd4543809536, 64'd301691168, - 64'd728253792256, - 64'd2209112576, 64'd4391622656, 64'd302338336, - 64'd726433529856, - 64'd5058731520, 64'd4236464640, 64'd302617536, - 64'd723208503296, - 64'd7827677696, 64'd4078595328, 64'd302531328, - 64'd718619738112, - 64'd10513341440, 64'd3918274816, 64'd302082976, - 64'd712709439488, - 64'd13113285632, 64'd3755764480, 64'd301276256, - 64'd705521123328, - 64'd15625242624, 64'd3591326208, 64'd300115520, - 64'd697099223040, - 64'd18047119360, 64'd3425220608, 64'd298605664, - 64'd687489286144, - 64'd20376993792, 64'd3257708288, 64'd296752064, - 64'd676737843200, - 64'd22613118976, 64'd3089048576, 64'd294560736, - 64'd664892080128, - 64'd24753920000, 64'd2919499520, 64'd292038048, - 64'd652000034816, - 64'd26798000128, 64'd2749316608, 64'd289190944, - 64'd638110400512, - 64'd28744130560, 64'd2578753536, 64'd286026784, - 64'd623272394752, - 64'd30591258624, 64'd2408060928, 64'd282553408, - 64'd607535759360, - 64'd32338505728, 64'd2237486336, 64'd278778976, - 64'd590950694912, - 64'd33985155072, 64'd2067274112, 64'd274712192, - 64'd573567467520, - 64'd35530665984, 64'd1897664256, 64'd270361984, - 64'd555436933120, - 64'd36974665728, 64'd1728892928, 64'd265737808, - 64'd536609783808, - 64'd38316945408, 64'd1561191680, 64'd260849328, - 64'd517136941056, - 64'd39557451776, 64'd1394787200, 64'd255706560, - 64'd497069260800, - 64'd40696303616, 64'd1229901184, 64'd250319824, - 64'd476457533440, - 64'd41733771264, 64'd1066749632, 64'd244699744, - 64'd455352320000, - 64'd42670284800, 64'd905542912, 64'd238857120, - 64'd433803984896, - 64'd43506413568, 64'd746485440, 64'd232803056, - 64'd411862532096, - 64'd44242890752, 64'd589775296, 64'd226548832, - 64'd389577572352, - 64'd44880584704, 64'd435604288, 64'd220105888, - 64'd366998224896, - 64'd45420507136, 64'd284157280, 64'd213485872, - 64'd344173150208, - 64'd45863813120, 64'd135612352, 64'd206700560, - 64'd321150320640, - 64'd46211780608, - 64'd9859543, 64'd199761840, - 64'd297977020416, - 64'd46465826816, - 64'd152094736, 64'd192681680, - 64'd274699894784, - 64'd46627483648, - 64'd290937024, 64'd185472160, - 64'd251364671488, - 64'd46698405888, - 64'd426237760, 64'd178145408, - 64'd228016308224, - 64'd46680375296, - 64'd557856064, 64'd170713552, - 64'd204698812416, - 64'd46575267840, - 64'd685658880, 64'd163188784, - 64'd181455224832, - 64'd46385074176, - 64'd809521088, 64'd155583232, - 64'd158327570432, - 64'd46111883264, - 64'd929325632, 64'd147909040, - 64'd135356817408, - 64'd45757886464, - 64'd1044963584, 64'd140178272, - 64'd112582778880, - 64'd45325357056, - 64'd1156334208, 64'd132402944, - 64'd90044153856, - 64'd44816658432, - 64'd1263344768, 64'd124594992, - 64'd67778412544, - 64'd44234235904, - 64'd1365911168, 64'd116766208, - 64'd45821788160, - 64'd43580604416, - 64'd1463957248, 64'd108928312, - 64'd24209246208, - 64'd42858356736, - 64'd1557415168, 64'd101092824, - 64'd2974428672, - 64'd42070142976, - 64'd1646225536, 64'd93271160, 64'd17850353664, - 64'd41218678784, - 64'd1730336896, 64'd85474520, 64'd38234165248, - 64'd40306724864, - 64'd1809705984, 64'd77713928, 64'd58147467264, - 64'd39337099264, - 64'd1884298112, 64'd70000208, 64'd77562126336, - 64'd38312656896, - 64'd1954086144, 64'd62343932, 64'd96451469312, - 64'd37236293632, - 64'd2019051008, 64'd54755468, 64'd114790252544, - 64'd36110934016, - 64'd2079181952, 64'd47244916, 64'd132554727424, - 64'd34939535360, - 64'd2134475520, 64'd39822112, 64'd149722611712, - 64'd33725071360, - 64'd2184935936, 64'd32496616, 64'd166273122304, - 64'd32470532096, - 64'd2230575616, 64'd25277704, 64'd182186967040, - 64'd31178921984, - 64'd2271413760, 64'd18174346, 64'd197446352896, - 64'd29853249536, - 64'd2307476992, 64'd11195207, 64'd212035026944, - 64'd28496527360, - 64'd2338799104, 64'd4348626, 64'd225938210816, - 64'd27111757824, - 64'd2365421056, - 64'd2357381, 64'd239142617088, - 64'd25701941248, - 64'd2387390208, - 64'd8915142, 64'd251636465664, - 64'd24270059520, - 64'd2404760576, - 64'd15317325, 64'd263409483776, - 64'd22819080192, - 64'd2417593088, - 64'd21556954, 64'd274452856832, - 64'd21351946240, - 64'd2425954048, - 64'd27627412, 64'd284759228416, - 64'd19871571968, - 64'd2429916672, - 64'd33522442, 64'd294322700288, - 64'd18380845056, - 64'd2429559296, - 64'd39236160, 64'd303138832384, - 64'd16882610176, - 64'd2424966144, - 64'd44763060, 64'd311204511744, - 64'd15379678208, - 64'd2416226560, - 64'd50098004, 64'd318518165504, - 64'd13874812928, - 64'd2403435264, - 64'd55236240, 64'd325079465984, - 64'd12370733056, - 64'd2386691840, - 64'd60173392, 64'd330889494528, - 64'd10870104064, - 64'd2366100224, - 64'd64905476, 64'd335950577664, - 64'd9375537152, - 64'd2341769216, - 64'd69428888, 64'd340266450944, - 64'd7889585664, - 64'd2313811200, - 64'd73740416, 64'd343842029568, - 64'd6414739968, - 64'd2282343168, - 64'd77837216, 64'd346683441152, - 64'd4953428480, - 64'd2247484928, - 64'd81716832, 64'd348798091264, - 64'd3508009728, - 64'd2209360640, - 64'd85377208, 64'd350194499584, - 64'd2080774016, - 64'd2168096512, - 64'd88816648, 64'd350882267136, - 64'd673937472, - 64'd2123822848, - 64'd92033824, 64'd350872174592, 64'd710358208, - 64'd2076671616, - 64'd95027808, 64'd350176018432, 64'd2070049152, - 64'd2026777600, - 64'd97798024, 64'd348806545408, 64'd3403151104, - 64'd1974277376, - 64'd100344256, 64'd346777616384, 64'd4707761152, - 64'd1919309952, - 64'd102666648, 64'd344103845888, 64'd5982059520, - 64'd1862015232, - 64'd104765704, 64'd340800897024, 64'd7224311808, - 64'd1802534912, - 64'd106642272, 64'd336885153792, 64'd8432869888, - 64'd1741011712, - 64'd108297536, 64'd332373884928, 64'd9606172672, - 64'd1677589120, - 64'd109733016, 64'd327285112832, 64'd10742748160, - 64'd1612411136, - 64'd110950552, 64'd321637482496, 64'd11841213440, - 64'd1545622144, - 64'd111952312, 64'd315450458112, 64'd12900276224, - 64'd1477366784, - 64'd112740760, 64'd308743995392, 64'd13918737408, - 64'd1407789440, - 64'd113318664, 64'd301538672640, 64'd14895484928, - 64'd1337033984, - 64'd113689088, 64'd293855625216, 64'd15829501952, - 64'd1265243904, - 64'd113855368, 64'd285716447232, 64'd16719862784, - 64'd1192561792, - 64'd113821120, 64'd277143191552, 64'd17565732864, - 64'd1119129088, - 64'd113590208, 64'd268158255104, 64'd18366367744, - 64'd1045086016, - 64'd113166760, 64'd258784460800, 64'd19121117184, - 64'd970571456, - 64'd112555144, 64'd249044877312, 64'd19829422080, - 64'd895722432, - 64'd111759944, 64'd238962851840, 64'd20490811392, - 64'd820674112, - 64'd110785976, 64'd228561944576, 64'd21104902144, - 64'd745559744, - 64'd109638248, 64'd217865879552, 64'd21671403520, - 64'd670510080, - 64'd108321976, 64'd206898511872, 64'd22190108672, - 64'd595653696, - 64'd106842552, 64'd195683762176, 64'd22660902912, - 64'd521116320, - 64'd105205544, 64'd184245600256, 64'd23083747328, - 64'd447021088, - 64'd103416680, 64'd172607995904, 64'd23458697216, - 64'd373488128, - 64'd101481824, 64'd160794869760, 64'd23785879552, - 64'd300634528, - 64'd99407000, 64'd148830044160, 64'd24065511424, - 64'd228574128, - 64'd97198328, 64'd136737234944, 64'd24297881600, - 64'd157417440, - 64'd94862056, 64'd124539977728, 64'd24483358720, - 64'd87271464, - 64'd92404536, 64'd112261619712, 64'd24622387200, - 64'd18239634, - 64'd89832192, 64'd99925254144, 64'd24715481088, 64'd49578332, - 64'd87151536, 64'd87553695744, 64'd24763226112, 64'd116086544, - 64'd84369136, 64'd75169472512, 64'd24766281728, 64'd181192992, - 64'd81491624, 64'd62794747904, 64'd24725364736, 64'd244809696, - 64'd78525664, 64'd50451308544, 64'd24641265664, 64'd306852736, - 64'd75477936, 64'd38160543744, 64'd24514826240, 64'd367242272, - 64'd72355168, 64'd25943390208, 64'd24346955776, 64'd425902784, - 64'd69164072, 64'd13820332032, 64'd24138616832, 64'd482762944, - 64'd65911356, 64'd1811350400, 64'd23890825216, 64'd537755776, - 64'd62603716, - 64'd10064093184, 64'd23604645888, 64'd590818496, - 64'd59247820, - 64'd21787082752, 64'd23281199104, 64'd641892992, - 64'd55850300, - 64'd33339271168, 64'd22921641984, 64'd690925248, - 64'd52417744, - 64'd44702904320, 64'd22527182848, 64'd737865792, - 64'd48956668, - 64'd55860842496, 64'd22099064832, 64'd782669696, - 64'd45473540, - 64'd66796572672, 64'd21638572032, 64'd825296256, - 64'd41974736, - 64'd77494239232, 64'd21147019264, 64'd865709248, - 64'd38466552, - 64'd87938637824, 64'd20625756160, 64'd903876928, - 64'd34955184, - 64'd98115272704, 64'd20076163072, 64'd939771840, - 64'd31446734, - 64'd108010307584, 64'd19499638784, 64'd973370944, - 64'd27947182, - 64'd117610659840, 64'd18897614848, 64'd1004655424, - 64'd24462388, - 64'd126903918592, 64'd18271537152, 64'd1033610880, - 64'd20998092, - 64'd135878426624, 64'd17622872064, 64'd1060227008, - 64'd17559890, - 64'd144523264000, 64'd16953097216, 64'd1084497792, - 64'd14153241, - 64'd152828248064, 64'd16263705600, 64'd1106421120, - 64'd10783452, - 64'd160783958016, 64'd15556200448, 64'd1125999232, - 64'd7455676, - 64'd168381677568, 64'd14832087040, 64'd1143238144, - 64'd4174906, - 64'd175613526016, 64'd14092879872, 64'd1158147712, - 64'd945966, - 64'd182472294400, 64'd13340089344, 64'd1170741760, 64'd2226493, - 64'd188951592960, 64'd12575229952, 64'd1181037824, 64'd5337993, - 64'd195045769216, 64'd11799806976, 64'd1189057024, 64'd8384241, - 64'd200749891584, 64'd11015324672, 64'd1194823808, 64'd11361127, - 64'd206059831296, 64'd10223272960, 64'd1198366464, 64'd14264733, - 64'd210972147712, 64'd9425134592, 64'd1199716352, 64'd17091330, - 64'd215484186624, 64'd8622377984, 64'd1198908160, 64'd19837388, - 64'd219593998336, 64'd7816452608, 64'd1195979520, 64'd22499570, - 64'd223300354048, 64'd7008794112, 64'd1190971136, 64'd25074746, - 64'd226602745856, 64'd6200815104, 64'd1183926656, 64'd27559984, - 64'd229501353984, 64'd5393906688, 64'd1174892416, 64'd29952556, - 64'd231997046784, 64'd4589435904, 64'd1163917312, 64'd32249940, - 64'd234091413504, 64'd3788742912, 64'd1151052928, 64'd34449816, - 64'd235786649600, 64'd2993140224, 64'd1136353024, 64'd36550072, - 64'd237085605888, 64'd2203910400, 64'd1119873664, 64'd38548808, - 64'd237991821312, 64'd1422304256, 64'd1101672960, 64'd40444320, - 64'd238509391872, 64'd649539328, 64'd1081811200, 64'd42235112, - 64'd238643036160, - 64'd113201360, 64'd1060350080, 64'd43919896, - 64'd238398046208, - 64'd864771136, 64'd1037353472, 64'd45497580, - 64'd237780303872, - 64'd1604060800, 64'd1012886464, 64'd46967280, - 64'd236796215296, - 64'd2329999872, 64'd987015808, 64'd48328308, - 64'd235452710912, - 64'd3041558016, 64'd959809408, 64'd49580176, - 64'd233757212672, - 64'd3737746176, 64'd931336320, 64'd50722580, - 64'd231717683200, - 64'd4417616896, 64'd901666624, 64'd51755424, - 64'd229342461952, - 64'd5080265728, 64'd870871360, 64'd52678784, - 64'd226640429056, - 64'd5724833280, 64'd839022144, 64'd53492940, - 64'd223620792320, - 64'd6350503424, 64'd806191424, 64'd54198332, - 64'd220293201920, - 64'd6956505600, 64'd772451904, 64'd54795596, - 64'd216667684864, - 64'd7542115840, 64'd737876800, 64'd55285532, - 64'd212754595840, - 64'd8106655744, 64'd702539392, 64'd55669116, - 64'd208564633600, - 64'd8649493504, 64'd666513216, 64'd55947480, - 64'd204108808192, - 64'd9170045952, 64'd629871616, 64'd56121928, - 64'd199398391808, - 64'd9667774464, 64'd592687872, 64'd56193908, - 64'd194444918784, - 64'd10142189568, 64'd555034944, 64'd56165024, - 64'd189260169216, - 64'd10592849920, 64'd516985344, 64'd56037028, - 64'd183856103424, - 64'd11019360256, 64'd478611136, 64'd55811808, - 64'd178244894720, - 64'd11421373440, 64'd439983712, 64'd55491384, - 64'd172438863872, - 64'd11798588416, 64'd401173696, 64'd55077908, - 64'd166450479104, - 64'd12150753280, 64'd362250944, 64'd54573656, - 64'd160292323328, - 64'd12477660160, 64'd323284256, 64'd53981016, - 64'd153977044992, - 64'd12779149312, 64'd284341408, 64'd53302488, - 64'd147517423616, - 64'd13055105024, 64'd245489072, 64'd52540680, - 64'd140926222336, - 64'd13305457664, 64'd206792592, 64'd51698296, - 64'd134216237056, - 64'd13530182656, 64'd168316000, 64'd50778136, - 64'd127400304640, - 64'd13729299456, 64'd130121920, 64'd49783076, - 64'd120491196416, - 64'd13902867456, 64'd92271440, 64'd48716084, - 64'd113501675520, - 64'd14050993152, 64'd54824076, 64'd47580192, - 64'd106444423168, - 64'd14173821952, 64'd17837676, 64'd46378508, - 64'd99332038656, - 64'd14271538176, - 64'd18631644, 64'd45114188, - 64'd92177031168, - 64'd14344369152, - 64'd54529576, 64'd43790452, - 64'd84991770624, - 64'd14392578048, - 64'd89803664, 64'd42410568, - 64'd77788504064, - 64'd14416467968, - 64'd124403384, 64'd40977836, - 64'd70579306496, - 64'd14416375808, - 64'd158280192, 64'd39495604, - 64'd63376064512, - 64'd14392675328, - 64'd191387552, 64'd37967240, - 64'd56190496768, - 64'd14345773056, - 64'd223681008, 64'd36396140, - 64'd49034088448, - 64'd14276109312, - 64'd255118208, 64'd34785712, - 64'd41918103552, - 64'd14184155136, - 64'd285658976, 64'd33139376, - 64'd34853564416, - 64'd14070413312, - 64'd315265312, 64'd31460558, - 64'd27851235328, - 64'd13935413248, - 64'd343901376, 64'd29752682, - 64'd20921602048, - 64'd13779713024, - 64'd371533664, 64'd28019164, - 64'd14074874880, - 64'd13603896320, - 64'd398130784, 64'd26263408, - 64'd7320958464, - 64'd13408571392, - 64'd423663776, 64'd24488800, - 64'd669450048, - 64'd13194371072, - 64'd448105888, 64'd22698702, 64'd5870374912, - 64'd12961948672, - 64'd471432608, 64'd20896444, 64'd12289572864, - 64'd12711977984, - 64'd493621792, 64'd19085330, 64'd18579542016, - 64'd12445151232, - 64'd514653600, 64'd17268614, 64'd24732033024, - 64'd12162180096, - 64'd534510400, 64'd15449513, 64'd30739152896, - 64'd11863788544, - 64'd553176960, 64'd13631193, 64'd36593373184, - 64'd11550717952, - 64'd570640256, 64'd11816766};
endpackage
`endif
