`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam N = 4;
	localparam real Lfr[0:3] = {[0.98584214], [0.98584214], [0.97811711], [0.97811711]};
	localparam real Lfi[0:3] = {[0.10665247], [-0.10665247], [0.04106261], [-0.04106261]};
	localparam real Lbr[0:3] = {[0.98584214], [0.98584214], [0.97811711], [0.97811711]};
	localparam real Lbi[0:3] = {[0.10665247], [-0.10665247], [0.04106261], [-0.04106261]};
	localparam real Wfr[0:3] = {[8.59515477e-05], [8.59515477e-05], [-2.80217754e-05], [-2.80217754e-05]};
	localparam real Wfi[0:3] = {[0.00010408], [-0.00010408], [-0.00011769], [0.00011769]};
	localparam real Wbr[0:3] = {[-8.59515477e-05], [-8.59515477e-05], [2.80217754e-05], [2.80217754e-05]};
	localparam real Wbi[0:3] = {[-0.00010408], [0.00010408], [0.00011769], [-0.00011769]};
	localparam real Ffr[0:3][0:79] = '{
		'{9.517403442589092, 5.803958733344014, -0.4775028600506327, -0.051475557707039, 12.334175399393775, 5.453185696094708, -0.5490632879926326, -0.04322707994592666, 14.96102263415146, 5.045163100567296, -0.6130702424751429, -0.03461632419982426, 17.37071831975333, 4.585572275315287, -0.6689092796911043, -0.025749026363305512, 19.53900499187631, 4.080596352735773, -0.7160707871752784, -0.01673212178091013, 21.444825625147537, 3.5368402976503113, -0.7541541277356487, -0.007672487370335698, 23.070513795269598, 2.9612473918572286, -0.7828704526032709, 0.0013242945205483789, 24.401941410865636, 2.3610132006917723, -0.8020441735158046, 0.010155136578104976, 25.428623015324696, 1.7434980596004206, -0.8116130991452264, 0.018720598010421204, 26.143776178374335, 1.1161391184899858, -0.8116272566501304, 0.02692597454909598, 26.544338013417295, 0.486362969358328, -0.802246434005084, 0.03468231537764404, 26.630938363918823, -0.1385001412055984, -0.7837364929699213, 0.04190735643865942, 26.407830694600133, -0.7512995481769507, -0.7564645159572013, 0.048526360716390216, 25.882782195429897, -1.345143932141644, -0.7208928624949469, 0.05447285732557144, 25.066925053280514, -1.913476746075026, -0.677572222336209, 0.05968927254545548, 23.974571262882375, -2.4501465043811197, -0.6271337624237217, 0.06412744730359313, 22.622993731046726, -2.949471206591621, -0.5702804737794054, 0.06774903702028089, 21.03217677218664, -3.406296248196691, -0.5077778318738266, 0.0705257911547416, 19.224539395604726, -3.8160452573072905, -0.4404438900763632, 0.07243971123109369, 17.224635043031086, -4.174763387130108, -0.36913893034683815, 0.0734830875492399},
		'{9.51740344258746, 5.803958733344131, -0.47750286005066395, -0.05147555770703265, 12.334175399392215, 5.45318569609482, -0.5490632879926624, -0.043227079945920587, 14.961022634149993, 5.045163100567405, -0.613070242475171, -0.03461632419981855, 17.37071831975197, 4.585572275315388, -0.6689092796911302, -0.0257490263633002, 19.53900499187507, 4.080596352735866, -0.716070787175302, -0.016732121780905287, 21.444825625146432, 3.5368402976503965, -0.7541541277356698, -0.0076724873703313615, 23.07051379526864, 2.961247391857304, -0.7828704526032892, 0.0013242945205521675, 24.401941410864822, 2.361013200691838, -0.8020441735158201, 0.010155136578108175, 25.428623015324046, 1.743498059600476, -0.8116130991452388, 0.018720598010423785, 26.143776178373848, 1.1161391184900298, -0.8116272566501396, 0.026925974549097925, 26.544338013416983, 0.4863629693583609, -0.8022464340050901, 0.03468231537764534, 26.63093836391867, -0.1385001412055773, -0.7837364929699241, 0.041907356438660066, 26.407830694600147, -0.7512995481769416, -0.7564645159572009, 0.04852636071639022, 25.882782195430078, -1.3451439321416463, -0.7208928624949434, 0.054472857325570806, 25.06692505328085, -1.9134767460750393, -0.6775722223362024, 0.05968927254545422, 23.974571262882865, -2.450146504381144, -0.6271337624237122, 0.0641274473035913, 22.62299373104736, -2.949471206591656, -0.5702804737793931, 0.06774903702027849, 21.032176772187412, -3.406296248196736, -0.507777831873812, 0.07052579115473867, 19.224539395605618, -3.8160452573073442, -0.44044389007634605, 0.07243971123109028, 17.224635043032087, -4.17476338713017, -0.3691389303468188, 0.07348308754923608},
		'{-9.313313592773765, -5.688953814066472, 0.40599510904134345, -0.19382811981932202, -12.087015729293103, -5.405857783345071, 0.3589502986526131, -0.18671439091601966, -14.719161330735629, -5.1228350901578645, 0.31308546179083796, -0.17949236217734052, -17.209940666047885, -4.8404954274546945, 0.2684508079689891, -0.17218217464535937, -19.559842146665797, -4.559421645725951, 0.22509179460033948, -0.16480332234289366, -21.769638866145826, -4.280169607798952, 0.18304922627424028, -0.1573746369854663, -23.840375083421378, -4.003268108103177, 0.14235935997530536, -0.14991427476315658, -25.77335268129348, -3.7292188538971804, 0.10305401577095727, -0.14243970513484921, -27.570117630503294, -3.4584965059201647, 0.0651606925002054, -0.13496770157542248, -29.23244648845956, -3.191548775908135, 0.0287026880051382, -0.1275143342146665, -30.762332960409537, -2.9287965783978374, -0.006300776544155451, -0.12009496430516839, -32.16197454955081, -2.6706342342314704, -0.039834428670685595, -0.11272424045505701, -33.43375932128638, -2.417429723170744, -0.07188681338676661, -0.10541609656034238, -34.58025280553011, -2.169524983030432, -0.10245015918354083, -0.09818375137062299, -35.60418505967578, -1.927236252748512, -0.13152024162071368, -0.09103970962115071, -36.508437913554964, -1.6908544568223671, -0.15909624491166258, -0.0839957646636417, -37.2960324164273, -1.4606456285578837, -0.18518062188698006, -0.07706300252778789, -37.9701165047758, -1.2368513696004657, -0.2097789527070889, -0.07025180734515825, -38.53395290842061, -1.0196893432437162, -0.23289980268185642, -0.06357186806706984, -38.990907311220546, -0.8093537990426116, -0.2545545795421773, -0.05703218640805522},
		'{-9.313313592769488, -5.688953814066671, 0.40599510904141745, -0.1938281198193366, -12.08701572928894, -5.405857783345265, 0.35895029865268496, -0.18671439091603384, -14.71916133073158, -5.122835090158053, 0.31308546179090785, -0.1794923621773543, -17.209940666043956, -4.8404954274548775, 0.2684508079690569, -0.17218217464537272, -19.559842146661993, -4.559421645726127, 0.22509179460040502, -0.1648033223429066, -21.769638866142145, -4.280169607799123, 0.18304922627430356, -0.15737463698547874, -23.84037508341783, -4.0032681081033425, 0.14235935997536636, -0.14991427476316863, -25.773352681290067, -3.729218853897339, 0.10305401577101594, -0.14243970513486076, -27.570117630500015, -3.4584965059203165, 0.06516069250026163, -0.13496770157543359, -29.232446488456414, -3.191548775908281, 0.0287026880051921, -0.12751433421467714, -30.76233296040653, -2.9287965783979777, -0.0063007765441039365, -0.12009496430517856, -32.161974549547935, -2.6706342342316036, -0.039834428670636524, -0.1127242404550667, -33.43375932128365, -2.41742972317087, -0.07188681338671998, -0.10541609656035161, -34.580252805527515, -2.169524983030552, -0.10245015918349654, -0.09818375137063172, -35.60418505967332, -1.9272362527486258, -0.13152024162067183, -0.09103970962115898, -36.50843791355265, -1.6908544568224744, -0.1590962449116232, -0.0839957646636495, -37.29603241642513, -1.4606456285579843, -0.1851806218869431, -0.0770630025277952, -37.97011650477375, -1.23685136960056, -0.2097789527070543, -0.0702518073451651, -38.5339529084187, -1.0196893432438041, -0.23289980268182417, -0.06357186806707624, -38.99090731121877, -0.8093537990426936, -0.25455457954214733, -0.05703218640806115}};
localparam real Ffi[0:3][0:79] = '{
	'{-27.674164915298654, 2.5184733274811264, 0.7343556810658382, -0.07050651561734925, -26.267303371139647, 3.101823664729105, 0.6730319166502996, -0.07499828955147023, -24.57994429148466, 3.639504198693084, 0.6049442691826638, -0.07854674905514027, -22.636314861901248, 4.12605570931263, 0.5309940973721856, -0.08112661160071676, -20.463203071189568, 4.556702195122724, 0.4521355305666279, -0.08272422960131473, -18.089604766013927, 4.927394718959295, 0.3693635411114507, -0.0833375536092401, -15.546351057642116, 5.234846103754052, 0.2837017436183584, -0.08297596187978651, -12.865720722547834, 5.476556229982367, 0.1961900669407216, -0.08165996051034236, -10.081042334625243, 5.650827799274608, 0.10787244368610588, -0.07942075979239319, -7.226290906310707, 5.756772541325502, 0.01978465946861291, -0.07629973375248889, -4.335683799492918, 5.794307952239594, -0.06705750012583211, -0.0723477710935723, -1.4432805958451844, 5.764144760575793, -0.15166967264393882, -0.06762452686766418, 1.4174085081242387, 5.667765421397218, -0.2331097869118613, -0.06219758520374837, 4.213801391108748, 5.507394037457768, -0.310488259713732, -0.05614154427142712, 6.914605614918611, 5.2859581992078155, -0.3829774142141183, -0.04953703537388402, 9.490159050556638, 5.007043320611547, -0.44982002413274885, -0.042469688627054455, 11.912745930888414, 4.674840124971845, -0.5103368994063947, -0.035029058091642695, 14.156885082907731, 4.294086003296922, -0.5639334415784055, -0.027307519478572413, 16.199587468981022, 3.8700010265739313, -0.6101051102832953, -0.01939915364627895, 18.02058056976475, 3.408219442116292, -0.6484417557795994, -0.011398629051431363},
	'{27.674164915299137, -2.518473327481149, -0.7343556810658288, 0.07050651561734744, 26.267303371140297, -3.10182366472914, -0.673031916650287, 0.07499828955146777, 24.579944291485468, -3.63950419869313, -0.6049442691826482, 0.07854674905513719, 22.6363148619022, -4.126055709312688, -0.5309940973721673, 0.0811266116007131, 20.463203071190655, -4.556702195122791, -0.45213553056660705, 0.08272422960131058, 18.08960476601513, -4.927394718959372, -0.36936354111142766, 0.08333755360923549, 15.546351057643417, -5.234846103754137, -0.2837017436183335, 0.08297596187978151, 12.86572072254922, -5.476556229982458, -0.19619006694069507, 0.08165996051033703, 10.081042334626694, -5.650827799274705, -0.10787244368607801, 0.07942075979238758, 7.226290906312207, -5.756772541325604, -0.019784659468584098, 0.07629973375248308, 4.335683799494449, -5.7943079522396985, 0.06705750012586148, 0.07234777109356638, 1.443280595846728, -5.7641447605759, 0.15166967264396847, 0.06762452686765819, -1.4174085081226995, -5.667765421397324, 0.2331097869118908, 0.06219758520374241, -4.213801391107234, -5.507394037457875, 0.310488259713761, 0.056141544271421234, -6.914605614917137, -5.28595819920792, 0.38297741421414655, 0.04953703537387829, -9.49015905055522, -5.0070433206116505, 0.44982002413277594, 0.04246968862704894, -11.912745930887068, -4.674840124971943, 0.5103368994064205, 0.035029058091637456, -14.156885082906472, -4.294086003297015, 0.5639334415784296, 0.02730751947856751, -16.199587468979864, -3.8700010265740183, 0.6101051102833174, 0.01939915364627442, -18.020580569763702, -3.408219442116372, 0.6484417557796194, 0.011398629051427259},
	'{72.51131969922037, -3.8625231707022207, 0.929323822626333, -0.06994708325861936, 70.5421336889876, -4.011603326911038, 0.9256587549077067, -0.07637552839346037, 68.50214369362797, -4.145796515909857, 0.9201421065661662, -0.082371192286889, 66.39871179008813, -4.265431518949687, 0.9128628483284804, -0.08793909836754918, 64.23903113887704, -4.370854958184794, 0.903910065718909, -0.0930849871807982, 62.03011743793533, -4.462429804040693, 0.8933727614134688, -0.09781527412782093, 59.77880111623674, -4.54053390928278, 0.8813396659957791, -0.10213700750176719, 57.49172025324865, -4.605558571848607, 0.8678990571746913, -0.10605782689940811, 55.1753142093852, -4.657907128358656, 0.8531385875030785, -0.10958592208272783, 52.83581795166512, -4.697993580074422, 0.8371451206171207, -0.11272999236079786, 50.479257057937836, -4.7262412529287605, 0.8200045759961625, -0.11549920655822801, 48.11144338226526, -4.743081493112122, 0.8018017822247844, -0.11790316363245998, 45.7379713633386, -4.748952399559536, 0.7826203387210673, -0.11995185399817505, 43.36421495717219, -4.7442975945474615, 0.7625424858782165, -0.1216556216131318, 40.99532517474419, -4.729565033476708, 0.7416489835506792, -0.12302512687584188, 38.63622820474926, -4.7052058547881135, 0.7200189978007006, -0.12407131038163734, 36.29162410118614, -4.67167327083134, 0.6977299958068675, -0.1248053575798879, 33.96598601512404, -4.6294215003843755, 0.6748576488226227, -0.12523866437139655, 31.66355994967266, -4.578904743402131, 0.6514757430599522, -0.1253828036813429, 29.388365016920893, -4.520576198457048, 0.6276560983614967, -0.12524949303956054},
	'{-72.51131969922082, 3.8625231707022434, -0.9293238226263425, 0.06994708325862117, -70.54213368898823, 4.011603326911068, -0.925658754907719, 0.07637552839346275, -68.50214369362877, 4.145796515909895, -0.9201421065661813, 0.08237119228689191, -66.39871179008907, 4.265431518949732, -0.912862848328498, 0.08793909836755259, -64.2390311388781, 4.370854958184845, -0.903910065718929, 0.09308498718080209, -62.03011743793654, 4.46242980404075, -0.8933727614134911, 0.09781527412782526, -59.778801116238064, 4.540533909282843, -0.8813396659958035, 0.10213700750177193, -57.491720253250094, 4.605558571848675, -0.8678990571747176, 0.10605782689941325, -55.175314209386755, 4.65790712835873, -0.8531385875031068, 0.10958592208273332, -52.83581795166677, 4.697993580074499, -0.8371451206171505, 0.1127299923608037, -50.47925705793958, 4.726241252928842, -0.8200045759961939, 0.11549920655823415, -48.11144338226708, 4.743081493112207, -0.8018017822248172, 0.11790316363246642, -45.737971363340506, 4.7489523995596254, -0.7826203387211014, 0.11995185399818173, -43.36421495717416, 4.744297594547554, -0.7625424858782519, 0.12165562161313871, -40.995325174746235, 4.729565033476804, -0.7416489835507156, 0.12302512687584899, -38.63622820475136, 4.705205854788212, -0.7200189978007379, 0.12407131038164465, -36.29162410118829, 4.671673270831441, -0.6977299958069055, 0.12480535757989536, -33.96598601512623, 4.6294215003844785, -0.6748576488226614, 0.12523866437140418, -31.663559949674887, 4.5789047434022345, -0.6514757430599915, 0.12538280368135063, -29.388365016923153, 4.520576198457154, -0.6276560983615366, 0.12524949303956834}};
	localparam real Fbr[0:3][0:79] = '{
		'{-9.517403442589092, 5.803958733344014, 0.4775028600506327, -0.051475557707039, -12.334175399393775, 5.453185696094708, 0.5490632879926326, -0.04322707994592666, -14.96102263415146, 5.045163100567296, 0.6130702424751429, -0.03461632419982426, -17.37071831975333, 4.585572275315287, 0.6689092796911043, -0.025749026363305512, -19.53900499187631, 4.080596352735773, 0.7160707871752784, -0.01673212178091013, -21.444825625147537, 3.5368402976503113, 0.7541541277356487, -0.007672487370335698, -23.070513795269598, 2.9612473918572286, 0.7828704526032709, 0.0013242945205483789, -24.401941410865636, 2.3610132006917723, 0.8020441735158046, 0.010155136578104976, -25.428623015324696, 1.7434980596004206, 0.8116130991452264, 0.018720598010421204, -26.143776178374335, 1.1161391184899858, 0.8116272566501304, 0.02692597454909598, -26.544338013417295, 0.486362969358328, 0.802246434005084, 0.03468231537764404, -26.630938363918823, -0.1385001412055984, 0.7837364929699213, 0.04190735643865942, -26.407830694600133, -0.7512995481769507, 0.7564645159572013, 0.048526360716390216, -25.882782195429897, -1.345143932141644, 0.7208928624949469, 0.05447285732557144, -25.066925053280514, -1.913476746075026, 0.677572222336209, 0.05968927254545548, -23.974571262882375, -2.4501465043811197, 0.6271337624237217, 0.06412744730359313, -22.622993731046726, -2.949471206591621, 0.5702804737794054, 0.06774903702028089, -21.03217677218664, -3.406296248196691, 0.5077778318738266, 0.0705257911547416, -19.224539395604726, -3.8160452573072905, 0.4404438900763632, 0.07243971123109369, -17.224635043031086, -4.174763387130108, 0.36913893034683815, 0.0734830875492399},
		'{-9.51740344258746, 5.803958733344131, 0.47750286005066395, -0.05147555770703265, -12.334175399392215, 5.45318569609482, 0.5490632879926624, -0.043227079945920587, -14.961022634149993, 5.045163100567405, 0.613070242475171, -0.03461632419981855, -17.37071831975197, 4.585572275315388, 0.6689092796911302, -0.0257490263633002, -19.53900499187507, 4.080596352735866, 0.716070787175302, -0.016732121780905287, -21.444825625146432, 3.5368402976503965, 0.7541541277356698, -0.0076724873703313615, -23.07051379526864, 2.961247391857304, 0.7828704526032892, 0.0013242945205521675, -24.401941410864822, 2.361013200691838, 0.8020441735158201, 0.010155136578108175, -25.428623015324046, 1.743498059600476, 0.8116130991452388, 0.018720598010423785, -26.143776178373848, 1.1161391184900298, 0.8116272566501396, 0.026925974549097925, -26.544338013416983, 0.4863629693583609, 0.8022464340050901, 0.03468231537764534, -26.63093836391867, -0.1385001412055773, 0.7837364929699241, 0.041907356438660066, -26.407830694600147, -0.7512995481769416, 0.7564645159572009, 0.04852636071639022, -25.882782195430078, -1.3451439321416463, 0.7208928624949434, 0.054472857325570806, -25.06692505328085, -1.9134767460750393, 0.6775722223362024, 0.05968927254545422, -23.974571262882865, -2.450146504381144, 0.6271337624237122, 0.0641274473035913, -22.62299373104736, -2.949471206591656, 0.5702804737793931, 0.06774903702027849, -21.032176772187412, -3.406296248196736, 0.507777831873812, 0.07052579115473867, -19.224539395605618, -3.8160452573073442, 0.44044389007634605, 0.07243971123109028, -17.224635043032087, -4.17476338713017, 0.3691389303468188, 0.07348308754923608},
		'{9.313313592773765, -5.688953814066472, -0.40599510904134345, -0.19382811981932202, 12.087015729293103, -5.405857783345071, -0.3589502986526131, -0.18671439091601966, 14.719161330735629, -5.1228350901578645, -0.31308546179083796, -0.17949236217734052, 17.209940666047885, -4.8404954274546945, -0.2684508079689891, -0.17218217464535937, 19.559842146665797, -4.559421645725951, -0.22509179460033948, -0.16480332234289366, 21.769638866145826, -4.280169607798952, -0.18304922627424028, -0.1573746369854663, 23.840375083421378, -4.003268108103177, -0.14235935997530536, -0.14991427476315658, 25.77335268129348, -3.7292188538971804, -0.10305401577095727, -0.14243970513484921, 27.570117630503294, -3.4584965059201647, -0.0651606925002054, -0.13496770157542248, 29.23244648845956, -3.191548775908135, -0.0287026880051382, -0.1275143342146665, 30.762332960409537, -2.9287965783978374, 0.006300776544155451, -0.12009496430516839, 32.16197454955081, -2.6706342342314704, 0.039834428670685595, -0.11272424045505701, 33.43375932128638, -2.417429723170744, 0.07188681338676661, -0.10541609656034238, 34.58025280553011, -2.169524983030432, 0.10245015918354083, -0.09818375137062299, 35.60418505967578, -1.927236252748512, 0.13152024162071368, -0.09103970962115071, 36.508437913554964, -1.6908544568223671, 0.15909624491166258, -0.0839957646636417, 37.2960324164273, -1.4606456285578837, 0.18518062188698006, -0.07706300252778789, 37.9701165047758, -1.2368513696004657, 0.2097789527070889, -0.07025180734515825, 38.53395290842061, -1.0196893432437162, 0.23289980268185642, -0.06357186806706984, 38.990907311220546, -0.8093537990426116, 0.2545545795421773, -0.05703218640805522},
		'{9.313313592769488, -5.688953814066671, -0.40599510904141745, -0.1938281198193366, 12.08701572928894, -5.405857783345265, -0.35895029865268496, -0.18671439091603384, 14.71916133073158, -5.122835090158053, -0.31308546179090785, -0.1794923621773543, 17.209940666043956, -4.8404954274548775, -0.2684508079690569, -0.17218217464537272, 19.559842146661993, -4.559421645726127, -0.22509179460040502, -0.1648033223429066, 21.769638866142145, -4.280169607799123, -0.18304922627430356, -0.15737463698547874, 23.84037508341783, -4.0032681081033425, -0.14235935997536636, -0.14991427476316863, 25.773352681290067, -3.729218853897339, -0.10305401577101594, -0.14243970513486076, 27.570117630500015, -3.4584965059203165, -0.06516069250026163, -0.13496770157543359, 29.232446488456414, -3.191548775908281, -0.0287026880051921, -0.12751433421467714, 30.76233296040653, -2.9287965783979777, 0.0063007765441039365, -0.12009496430517856, 32.161974549547935, -2.6706342342316036, 0.039834428670636524, -0.1127242404550667, 33.43375932128365, -2.41742972317087, 0.07188681338671998, -0.10541609656035161, 34.580252805527515, -2.169524983030552, 0.10245015918349654, -0.09818375137063172, 35.60418505967332, -1.9272362527486258, 0.13152024162067183, -0.09103970962115898, 36.50843791355265, -1.6908544568224744, 0.1590962449116232, -0.0839957646636495, 37.29603241642513, -1.4606456285579843, 0.1851806218869431, -0.0770630025277952, 37.97011650477375, -1.23685136960056, 0.2097789527070543, -0.0702518073451651, 38.5339529084187, -1.0196893432438041, 0.23289980268182417, -0.06357186806707624, 38.99090731121877, -0.8093537990426936, 0.25455457954214733, -0.05703218640806115}};
localparam real Fbi[0:3][0:79] = '{
	'{27.674164915298654, 2.5184733274811264, -0.7343556810658382, -0.07050651561734925, 26.267303371139647, 3.101823664729105, -0.6730319166502996, -0.07499828955147023, 24.57994429148466, 3.639504198693084, -0.6049442691826638, -0.07854674905514027, 22.636314861901248, 4.12605570931263, -0.5309940973721856, -0.08112661160071676, 20.463203071189568, 4.556702195122724, -0.4521355305666279, -0.08272422960131473, 18.089604766013927, 4.927394718959295, -0.3693635411114507, -0.0833375536092401, 15.546351057642116, 5.234846103754052, -0.2837017436183584, -0.08297596187978651, 12.865720722547834, 5.476556229982367, -0.1961900669407216, -0.08165996051034236, 10.081042334625243, 5.650827799274608, -0.10787244368610588, -0.07942075979239319, 7.226290906310707, 5.756772541325502, -0.01978465946861291, -0.07629973375248889, 4.335683799492918, 5.794307952239594, 0.06705750012583211, -0.0723477710935723, 1.4432805958451844, 5.764144760575793, 0.15166967264393882, -0.06762452686766418, -1.4174085081242387, 5.667765421397218, 0.2331097869118613, -0.06219758520374837, -4.213801391108748, 5.507394037457768, 0.310488259713732, -0.05614154427142712, -6.914605614918611, 5.2859581992078155, 0.3829774142141183, -0.04953703537388402, -9.490159050556638, 5.007043320611547, 0.44982002413274885, -0.042469688627054455, -11.912745930888414, 4.674840124971845, 0.5103368994063947, -0.035029058091642695, -14.156885082907731, 4.294086003296922, 0.5639334415784055, -0.027307519478572413, -16.199587468981022, 3.8700010265739313, 0.6101051102832953, -0.01939915364627895, -18.02058056976475, 3.408219442116292, 0.6484417557795994, -0.011398629051431363},
	'{-27.674164915299137, -2.518473327481149, 0.7343556810658288, 0.07050651561734744, -26.267303371140297, -3.10182366472914, 0.673031916650287, 0.07499828955146777, -24.579944291485468, -3.63950419869313, 0.6049442691826482, 0.07854674905513719, -22.6363148619022, -4.126055709312688, 0.5309940973721673, 0.0811266116007131, -20.463203071190655, -4.556702195122791, 0.45213553056660705, 0.08272422960131058, -18.08960476601513, -4.927394718959372, 0.36936354111142766, 0.08333755360923549, -15.546351057643417, -5.234846103754137, 0.2837017436183335, 0.08297596187978151, -12.86572072254922, -5.476556229982458, 0.19619006694069507, 0.08165996051033703, -10.081042334626694, -5.650827799274705, 0.10787244368607801, 0.07942075979238758, -7.226290906312207, -5.756772541325604, 0.019784659468584098, 0.07629973375248308, -4.335683799494449, -5.7943079522396985, -0.06705750012586148, 0.07234777109356638, -1.443280595846728, -5.7641447605759, -0.15166967264396847, 0.06762452686765819, 1.4174085081226995, -5.667765421397324, -0.2331097869118908, 0.06219758520374241, 4.213801391107234, -5.507394037457875, -0.310488259713761, 0.056141544271421234, 6.914605614917137, -5.28595819920792, -0.38297741421414655, 0.04953703537387829, 9.49015905055522, -5.0070433206116505, -0.44982002413277594, 0.04246968862704894, 11.912745930887068, -4.674840124971943, -0.5103368994064205, 0.035029058091637456, 14.156885082906472, -4.294086003297015, -0.5639334415784296, 0.02730751947856751, 16.199587468979864, -3.8700010265740183, -0.6101051102833174, 0.01939915364627442, 18.020580569763702, -3.408219442116372, -0.6484417557796194, 0.011398629051427259},
	'{-72.51131969922037, -3.8625231707022207, -0.929323822626333, -0.06994708325861936, -70.5421336889876, -4.011603326911038, -0.9256587549077067, -0.07637552839346037, -68.50214369362797, -4.145796515909857, -0.9201421065661662, -0.082371192286889, -66.39871179008813, -4.265431518949687, -0.9128628483284804, -0.08793909836754918, -64.23903113887704, -4.370854958184794, -0.903910065718909, -0.0930849871807982, -62.03011743793533, -4.462429804040693, -0.8933727614134688, -0.09781527412782093, -59.77880111623674, -4.54053390928278, -0.8813396659957791, -0.10213700750176719, -57.49172025324865, -4.605558571848607, -0.8678990571746913, -0.10605782689940811, -55.1753142093852, -4.657907128358656, -0.8531385875030785, -0.10958592208272783, -52.83581795166512, -4.697993580074422, -0.8371451206171207, -0.11272999236079786, -50.479257057937836, -4.7262412529287605, -0.8200045759961625, -0.11549920655822801, -48.11144338226526, -4.743081493112122, -0.8018017822247844, -0.11790316363245998, -45.7379713633386, -4.748952399559536, -0.7826203387210673, -0.11995185399817505, -43.36421495717219, -4.7442975945474615, -0.7625424858782165, -0.1216556216131318, -40.99532517474419, -4.729565033476708, -0.7416489835506792, -0.12302512687584188, -38.63622820474926, -4.7052058547881135, -0.7200189978007006, -0.12407131038163734, -36.29162410118614, -4.67167327083134, -0.6977299958068675, -0.1248053575798879, -33.96598601512404, -4.6294215003843755, -0.6748576488226227, -0.12523866437139655, -31.66355994967266, -4.578904743402131, -0.6514757430599522, -0.1253828036813429, -29.388365016920893, -4.520576198457048, -0.6276560983614967, -0.12524949303956054},
	'{72.51131969922082, 3.8625231707022434, 0.9293238226263425, 0.06994708325862117, 70.54213368898823, 4.011603326911068, 0.925658754907719, 0.07637552839346275, 68.50214369362877, 4.145796515909895, 0.9201421065661813, 0.08237119228689191, 66.39871179008907, 4.265431518949732, 0.912862848328498, 0.08793909836755259, 64.2390311388781, 4.370854958184845, 0.903910065718929, 0.09308498718080209, 62.03011743793654, 4.46242980404075, 0.8933727614134911, 0.09781527412782526, 59.778801116238064, 4.540533909282843, 0.8813396659958035, 0.10213700750177193, 57.491720253250094, 4.605558571848675, 0.8678990571747176, 0.10605782689941325, 55.175314209386755, 4.65790712835873, 0.8531385875031068, 0.10958592208273332, 52.83581795166677, 4.697993580074499, 0.8371451206171505, 0.1127299923608037, 50.47925705793958, 4.726241252928842, 0.8200045759961939, 0.11549920655823415, 48.11144338226708, 4.743081493112207, 0.8018017822248172, 0.11790316363246642, 45.737971363340506, 4.7489523995596254, 0.7826203387211014, 0.11995185399818173, 43.36421495717416, 4.744297594547554, 0.7625424858782519, 0.12165562161313871, 40.995325174746235, 4.729565033476804, 0.7416489835507156, 0.12302512687584899, 38.63622820475136, 4.705205854788212, 0.7200189978007379, 0.12407131038164465, 36.29162410118829, 4.671673270831441, 0.6977299958069055, 0.12480535757989536, 33.96598601512623, 4.6294215003844785, 0.6748576488226614, 0.12523866437140418, 31.663559949674887, 4.5789047434022345, 0.6514757430599915, 0.12538280368135063, 29.388365016923153, 4.520576198457154, 0.6276560983615366, 0.12524949303956834}};
	localparam real hf[0:3999] = {0.024986578, -0.000116877105, -3.896343e-05, 2.2712003e-07, 0.024869869, -0.0003495672, -3.6725352e-05, 6.683011e-07, 0.02463752, -0.00057908345, -3.2282736e-05, 1.071189e-06, 0.02429164, -0.00080335606, -2.5699466e-05, 1.4122909e-06, 0.023835355, -0.0010203768, -1.7068134e-05, 1.6701244e-06, 0.023272775, -0.0012282217, -6.508329e-06, 1.825436e-06, 0.02260895, -0.0014250721, 5.835373e-06, 1.8613864e-06, 0.021849804, -0.0016092348, 1.979567e-05, 1.7637041e-06, 0.021002075, -0.0017791594, 3.5185032e-05, 1.5208042e-06, 0.020073237, -0.0019334549, 5.1798383e-05, 1.1238726e-06, 0.019071415, -0.0020709035, 6.941594e-05, 5.669145e-07, 0.018005302, -0.0021904726, 8.7806206e-05, -1.5323168e-07, 0.016884053, -0.0022913238, 0.000106729, -1.0369153e-06, 0.015717195, -0.0023728213, 0.00012593858, -2.0817276e-06, 0.014514523, -0.0024345345, 0.00014518676, -3.2825897e-06, 0.01328599, -0.0024762424, 0.000164226, -4.6318687e-06, 0.012041612, -0.0024979326, 0.00018281244, -6.119525e-06, 0.010791358, -0.0024997983, 0.00020070883, -7.733287e-06, 0.009545049, -0.0024822343, 0.00021768737, -9.458844e-06, 0.008312262, -0.0024458296, 0.00023353235, -1.1280068e-05, 0.0071022296, -0.0023913574, 0.00024804258, -1.31792485e-05, 0.0059237573, -0.0023197657, 0.0002610337, -1.5137347e-05, 0.004785133, -0.0022321627, 0.00027234023, -1.7134254e-05, 0.003694055, -0.002129803, 0.00028181716, -1.9149073e-05, 0.0026575602, -0.0020140712, 0.0002893417, -2.116038e-05, 0.0016819648, -0.0018864649, 0.00029481426, -2.3146522e-05, 0.0007728115, -0.0017485761, 0.00029815955, -2.5085883e-05, -6.517271e-05, -0.0016020724, 0.00029932705, -2.6957157e-05, -0.0008281093, -0.0014486772, 0.0002982914, -2.8739623e-05, -0.0015129913, -0.0012901495, 0.00029505236, -3.0413386e-05, -0.002117696, -0.0011282647, 0.0002896347, -3.195963e-05, -0.0026409882, -0.00096479343, 0.0002820874, -3.3360822e-05, -0.003082513, -0.00080148317, 0.00027248287, -3.4600955e-05, -0.0034427792, -0.00064003846, 0.000260916, -3.5665686e-05, -0.0037231334, -0.0004821034, 0.00024750258, -3.6542533e-05, -0.003925726, -0.00032924407, 0.00023237792, -3.7221005e-05, -0.004053466, -0.00018293266, 0.00021569492, -3.76927e-05, -0.0041099745, -4.453296e-05, 0.00019762217, -3.79514e-05, -0.0040995227, 8.471297e-05, 0.00017834186, -3.7993144e-05, -0.0040269704, 0.00020369625, 0.00015804752, -3.7816237e-05, -0.0038976963, 0.00031145103, 0.00013694167, -3.742127e-05, -0.0037175252, 0.00040716256, 0.00011523339, -3.6811085e-05, -0.0034926496, 0.0004901733, 9.3135954e-05, -3.599074e-05, -0.0032295508, 0.00055998715, 7.086427e-05, -3.4967423e-05, -0.002934917, 0.0006162719, 4.8632493e-05, -3.3750366e-05, -0.0026155617, 0.0006588598, 2.6651622e-05, -3.235072e-05, -0.0022783414, 0.0006877456, 5.1271536e-06, -3.0781408e-05, -0.0019300748, 0.00070308376, -1.5743133e-05, -2.9056979e-05, -0.0015774649, 0.0007051833, -3.577129e-05, -2.7193415e-05, -0.0012270228, 0.00069450086, -5.4781158e-05, -2.5207955e-05, -0.00088499615, 0.00067163265, -7.261017e-05, -2.311889e-05, -0.00055730145, 0.0006373044, -8.911096e-05, -2.0945343e-05, -0.0002494623, 0.00059236056, -0.00010415277, -1.8707058e-05, 3.3447053e-05, 0.00053775206, -0.00011762269, -1.6424181e-05, 0.00028685166, 0.00047452268, -0.00012942658, -1.4117025e-05, 0.0005067189, 0.00040379557, -0.0001394899, -1.1805854e-05, 0.00068959437, 0.00032675808, -0.00014775814, -9.510665e-06, 0.0008326304, 0.00024464677, -0.00015419716, -7.2509692e-06, 0.0009336064, 0.00015873181, -0.00015879319, -5.0455933e-06, 0.0009909424, 7.03015e-05, -0.0001615527, -2.9124817e-06, 0.0010037036, -1.9353303e-05, -0.00016250192, -8.6851696e-07, 0.000971598, -0.00010895448, -0.00016168621, 1.0706473e-06, 0.00089496677, -0.00019725144, -0.00015916926, 2.890736e-06, 0.0007747661, -0.0002830354, -0.00015503199, 4.578985e-06, 0.0006125435, -0.0003651528, -0.0001493714, 6.1242554e-06, 0.00041040673, -0.00044251818, -0.00014229909, 7.517124e-06, 0.00017098685, -0.0005141254, -0.00013393987, 8.749958e-06, -0.000102604055, -0.0005790583, -0.00012442996, 9.816967e-06, -0.00040682033, -0.00063650013, -0.00011391535, 1.0714228e-05, -0.0007377343, -0.00068574096, -0.000102549915, 1.1439698e-05, -0.0010910918, -0.00072618475, -9.049353e-05, 1.1993197e-05, -0.0014623696, -0.0007573539, -7.791015e-05, 1.237638e-05, -0.0018468365, -0.0007788933, -6.496585e-05, 1.2592673e-05, -0.002239615, -0.0007905721, -5.1826923e-05, 1.2647208e-05, -0.0026357428, -0.0007922844, -3.8657945e-05, 1.2546729e-05, -0.0030302363, -0.00078404846, -2.5619947e-05, 1.22994825e-05, -0.0034181513, -0.0007660045, -1.2868641e-05, 1.1915097e-05, -0.0037946438, -0.0007384107, -5.527264e-07, 1.1404446e-05, -0.0041550267, -0.00070163846, 1.1187671e-05, 1.0779499e-05, -0.0044948263, -0.000656166, 2.2222448e-05, 1.0053163e-05, -0.004809833, -0.00060257106, 3.2432832e-05, 9.239121e-06, -0.005096149, -0.0005415224, 4.1712527e-05, 8.351654e-06, -0.0053502326, -0.00047377063, 4.9968694e-05, 7.4054738e-06, -0.0055689337, -0.0004001377, 5.7122783e-05, 6.415538e-06, -0.005749531, -0.00032150644, 6.311115e-05, 5.3968797e-06, -0.005889757, -0.00023880896, 6.788551e-05, 4.3644327e-06, -0.005987819, -0.00015301503, 7.1413204e-05, 3.33286e-06, -0.0060424167, -6.5120075e-05, 7.367729e-05, 2.3163923e-06, -0.0060527516, 2.3866987e-05, 7.467643e-05, 1.3286729e-06, -0.006018531, 0.00011293571, 7.442458e-05, 3.8261123e-07, -0.0059399647, 0.00020108608, 7.295059e-05, -5.097503e-07, -0.005817757, 0.00028734, 7.029756e-05, -1.3373586e-06, -0.0056530945, 0.00037075247, 6.652203e-05, -2.0902578e-06, -0.005447625, 0.00045042214, 6.169313e-05, -2.759682e-06, -0.0052034347, 0.00052550115, 5.589148e-05, -3.3381343e-06, -0.004923017, 0.00059520424, 4.9208058e-05, -3.819447e-06, -0.004609243, 0.00065881707, 4.1742933e-05, -4.198827e-06, -0.0042653196, 0.0007157032, 3.3603916e-05, -4.472884e-06, -0.003894752, 0.0007653107, 2.4905143e-05, -4.639643e-06, -0.0035012984, 0.0008071772, 1.5765636e-05, -4.698537e-06, -0.003088926, 0.0008409337, 6.307793e-06, -4.6503856e-06, -0.0026617618, 0.0008663077, -3.3441117e-06, -4.4973604e-06, -0.0022240446, 0.00088312494, -1.3065424e-05, -4.2429283e-06, -0.0017800763, 0.0008913099, -2.2732595e-05, -3.8917874e-06, -0.0013341709, 0.000890885, -3.2224616e-05, -3.4497868e-06, -0.0008906079, 0.00088196935, -4.142441e-05, -2.9238345e-06, -0.0004535831, 0.00086477544, -5.0220144e-05, -2.321794e-06, -2.7163756e-05, 0.00083960575, -5.850646e-05, -1.652374e-06, 0.00038475564, 0.0008068475, -6.618562e-05, -9.250065e-07, 0.0007784943, 0.0007669673, -7.316853e-05, -1.497222e-07, 0.0011506232, 0.00072050426, -7.937563e-05, 6.629815e-07, 0.0014979994, 0.000668063, -8.473774e-05, 1.5022744e-06, 0.0018177973, 0.0006103056, -8.919661e-05, 2.3571292e-06, 0.0021075346, 0.000547943, -9.270552e-05, 3.2164576e-06, 0.002365095, 0.00048172637, -9.522962e-05, 4.069244e-06, 0.002588746, 0.00041243774, -9.674611e-05, 4.9046766e-06, 0.0027771518, 0.00034088065, -9.7244396e-05, 5.7122747e-06, 0.0029293816, 0.00026787055, -9.672597e-05, 6.482007e-06, 0.0030449138, 0.00019422543, -9.520421e-05, 7.204406e-06, 0.0031236338, 0.00012075634, -9.270407e-05, 7.870673e-06, 0.0031658295, 4.8258335e-05, -8.926157e-05, 8.472772e-06, 0.0031721801, -2.2498389e-05, -8.492326e-05, 9.003513e-06, 0.003143742, -9.077683e-05, -7.974546e-05, 9.4566285e-06, 0.0030819303, -0.00015588106, -7.379349e-05, 9.826832e-06, 0.0029884963, -0.00021716346, -6.714076e-05, 1.0109866e-05, 0.0028655012, -0.00027403128, -5.9867805e-05, 1.030254e-05, 0.0027152882, -0.00032595254, -5.206122e-05, 1.0402753e-05, 0.0025404498, -0.000372461, -4.3812594e-05, 1.04095e-05, 0.0023437948, -0.0004131604, -3.5217337e-05, 1.032287e-05, 0.0021283112, -0.0004477277, -2.6373558e-05, 1.0144035e-05, 0.0018971302, -0.0004759157, -1.738085e-05, 9.875211e-06, 0.0016534871, -0.0004975543, -8.339134e-06, 9.5196265e-06, 0.001400683, -0.0005125514, 6.5249236e-07, 9.081469e-06, 0.0011420455, -0.00052089227, 9.4969e-06, 8.565822e-06, 0.00088089047, -0.00052263855, 1.810001e-05, 7.978593e-06, 0.00062048424, -0.0005179262, 2.6371838e-05, 7.3264337e-06, 0.00036400717, -0.0005069625, 3.422745e-05, 6.6166567e-06, 0.00011451893, -0.00049002253, 4.1587886e-05, 5.8571363e-06, -0.0001250745, -0.0004674449, 4.8380953e-05, 5.0562144e-06, -0.0003520511, -0.00043962628, 5.4541957e-05, 4.222595e-06, -0.0005639008, -0.00040701643, 6.0014332e-05, 3.365242e-06, -0.00075835024, -0.0003701115, 6.475016e-05, 2.4932692e-06, -0.0009333844, -0.00032944788, 6.871057e-05, 1.6158366e-06, -0.0010872651, -0.00028559507, 7.186606e-05, 7.4204394e-07, -0.0012185457, -0.00023914858, 7.419667e-05, -1.1917229e-07, -0.0013260824, -0.00019072261, 7.5692085e-05, -9.591386e-07, -0.0014090413, -0.00014094257, 7.635154e-05, -1.7695393e-06, -0.0014669029, -9.043767e-05, 7.6183744e-05, -2.5425059e-06, -0.0014994614, -3.9833558e-05, 7.5206575e-05, -3.2706998e-06, -0.0015068215, 1.0254878e-05, 7.344675e-05, -3.9473884e-06, -0.0014893912, 5.9230428e-05, 7.093935e-05, -4.566511e-06, -0.0014478713, 0.00010652019, 6.772732e-05, -5.122739e-06, -0.0013832418, 0.00015158176, 6.386082e-05, -5.6115227e-06, -0.0012967449, 0.00019390904, 5.93965e-05, -6.0291327e-06, -0.0011898658, 0.00023303744, 5.4396824e-05, -6.372689e-06, -0.0010643104, 0.00026854855, 4.8929178e-05, -6.6401776e-06, -0.0009219817, 0.0003000742, 4.3065043e-05, -6.830463e-06, -0.0007649533, 0.00032729987, 3.6879126e-05, -6.943284e-06, -0.00059544214, 0.00034996742, 3.0448418e-05, -6.9792427e-06, -0.00041577968, 0.00036787707, 2.3851286e-05, -6.9397847e-06, -0.0002283824, 0.00038088873, 1.716655e-05, -6.827166e-06, -3.5721743e-05, 0.0003889226, 1.0472569e-05, -6.6444177e-06, 0.00015970602, 0.00039195913, 3.84635e-06, -6.3952925e-06, 0.0003554097, 0.00039003804, -2.637314e-06, -6.0842167e-06, 0.0005489325, 0.000383257, -8.906665e-06, -5.7162215e-06, 0.0007378806, 0.00037176942, -1.4893752e-05, -5.2968808e-06, 0.00091995014, 0.0003557817, -2.0535148e-05, -4.8322336e-06, 0.0010929531, 0.00033554994, -2.5772597e-05, -4.328711e-06, 0.0012548412, 0.00031137612, -3.0553598e-05, -3.7930529e-06, 0.0014037276, 0.00028360382, -3.483191e-05, -3.2322278e-06, 0.0015379067, 0.00025261342, -3.8567974e-05, -2.653347e-06, 0.0016558714, 0.00021881713, -4.172925e-05, -2.0635835e-06, 0.0017563275, 0.00018265363, -4.4290467e-05, -1.4700853e-06, 0.0018382053, 0.0001445825, -4.6233796e-05, -8.798973e-07, 0.0019006693, 0.00010507852, -4.7548918e-05, -2.9988044e-07, 0.001943124, 6.462584e-05, -4.8233018e-05, 2.63363e-07, 0.0019652168, 2.3712253e-05, -4.829067e-05, 8.035608e-07, 0.001966839, -1.7176591e-05, -4.7733673e-05, 1.3148367e-06, 0.0019481225, -5.7562815e-05, -4.6580783e-05, 1.7917708e-06, 0.001909436, -9.6981734e-05, -4.4857356e-05, 2.229454e-06, 0.0018513753, -0.00013498706, -4.2594966e-05, 2.6235343e-06, 0.0017747541, -0.00017115581, -3.983091e-05, 2.9702587e-06, 0.0016805907, -0.00020509283, -3.6607682e-05, 3.2665032e-06, 0.0015700932, -0.00023643493, -3.2972388e-05, 3.5097996e-06, 0.0014446424, -0.00026485464, -2.8976121e-05, 3.6983504e-06, 0.0013057735, -0.00029006338, -2.4673294e-05, 3.8310386e-06, 0.0011551554, -0.0003118142, -2.012095e-05, 3.907428e-06, 0.0009945696, -0.00032990403, -1.537806e-05, 3.9277547e-06, 0.00082588807, -0.00034417518, -1.0504799e-05, 3.892914e-06, 0.0006510498, -0.0003545167, -5.5618216e-06, 3.8044357e-06, 0.00047203756, -0.0003608646, -6.095561e-07, 3.6644583e-06, 0.0002908543, -0.0003632021, 4.2925003e-06, 3.4756895e-06, 0.00010949978, -0.0003615589, 9.086454e-06, 3.2413664e-06, -7.005265e-05, -0.00035601013, 1.3716667e-05, 2.9652074e-06, -0.00024587815, -0.00034667485, 1.8130359e-05, 2.6513612e-06, -0.000416122, -0.00033371375, 2.2278178e-05, 2.3043497e-06, -0.00057901966, -0.00031732683, 2.6114716e-05, 1.929009e-06, -0.0007329159, -0.00029775038, 2.959897e-05, 1.5304275e-06, -0.00087628193, -0.00027525355, 3.269475e-05, 1.1138819e-06, -0.0010077311, -0.00025013494, 3.5371e-05, 6.847718e-07, -0.0011260324, -0.00022271842, 3.760211e-05, 2.4855487e-07, -0.0012301225, -0.00019334916, 3.936808e-05, -1.893183e-07, -0.001319115, -0.00016238925, 4.0654697e-05, -6.234677e-07, -0.0013923077, -0.0001302132, 4.1453575e-05, -1.0486458e-06, -0.0014491879, -9.720347e-05, 4.1762174e-05, -1.4597965e-06, -0.0014894352, -6.374589e-05, 4.1583724e-05, -1.8521115e-06, -0.0015129221, -3.0225176e-05, 4.092709e-05, -2.221082e-06, -0.0015197119, 2.9794865e-06, 3.980659e-05, -2.5625463e-06, -0.0015100557, 3.5498742e-05, 3.8241713e-05, -2.8727338e-06, -0.0014843857, 6.697716e-05, 3.6256835e-05, -3.1483007e-06, -0.0014433075, 9.707708e-05, 3.388084e-05, -3.386364e-06, -0.0013875904, 0.00012548224, 3.1146705e-05, -3.584526e-06, -0.0013181557, 0.00015190107, 2.8091063e-05, -3.740896e-06, -0.0012360639, 0.00017606962, 2.4753714e-05, -3.854103e-06, -0.0011424997, 0.00019775413, 2.1177106e-05, -3.9233023e-06, -0.0010387572, 0.00021675328, 1.74058e-05, -3.9481793e-06, -0.0009262218, 0.00023289995, 1.3485926e-05, -3.928943e-06, -0.0008063545, 0.00024606255, 9.464609e-06, -3.866315e-06, -0.0006806726, 0.00025614596, 5.3894196e-06, -3.7615139e-06, -0.0005507317, 0.00026309196, 1.3078055e-06, -3.6162312e-06, -0.00041810746, 0.00026687945, -2.7334515e-06, -3.4326067e-06, -0.00028437664, 0.00026752386, -6.688769e-06, -3.2131943e-06, -0.00015109948, 0.0002650765, -1.0514272e-05, -2.9609264e-06, -1.9801768e-05, 0.00025962334, -1.4168271e-05, -2.6790735e-06, 0.00010804198, 0.00025128332, -1.7611716e-05, -2.3712018e-06, 0.00023102465, 0.00024020665, -2.0808595e-05, -2.041126e-06, 0.0003478215, 0.00022657229, -2.3726312e-05, -1.6928611e-06, 0.000457204, 0.0002105856, -2.6336e-05, -1.3305736e-06, 0.00055805227, 0.0001924754, -2.86128e-05, -9.585298e-07, 0.0006493661, 0.00017249103, -3.053608e-05, -5.8104513e-07, 0.0007302744, 0.00015089898, -3.2089603e-05, -2.0243363e-07, 0.00080004294, 0.0001279797, -3.3261647e-05, 1.7304232e-07, 0.00085808046, 0.00010402399, -3.4045068e-05, 5.412203e-07, 0.000903943, 7.932951e-05, -3.4437293e-05, 8.9808447e-07, 0.0009373362, 5.4197226e-05, -3.4440294e-05, 1.2398096e-06, 0.00095811655, 2.8927887e-05, -3.4060486e-05, 1.5628023e-06, 0.00096629, 3.8185226e-06, -3.3308566e-05, 1.8637385e-06, 0.0009620094, -2.0840904e-05, -3.219934e-05, 2.139598e-06, 0.0009455702, -4.477073e-05, -3.075146e-05, 2.3876942e-06, 0.0009174042, -6.770467e-05, -2.8987177e-05, 2.6056998e-06, 0.00087807275, -8.939263e-05, -2.6931988e-05, 2.7916674e-06, 0.00082825747, -0.00010960339, -2.461432e-05, 2.9440466e-06, 0.0007687504, -0.00012812686, -2.2065136e-05, 3.0616948e-06, 0.0007004428, -0.00014477625, -1.9317536e-05, 3.1438838e-06, 0.0006243134, -0.00015938978, -1.6406348e-05, 3.1903023e-06, 0.000541415, -0.00017183211, -1.33676895e-05, 3.2010514e-06, 0.0004528613, -0.00018199554, -1.0238536e-05, 3.1766376e-06, 0.00035981278, -0.00018980069, -7.0562724e-06, 3.1179597e-06, 0.00026346243, -0.00019519699, -3.8582616e-06, 3.0262931e-06, 0.00016502131, -0.00019816274, -6.8140974e-07, 2.9032674e-06, 6.570411e-05, -0.00019870495, 2.4382505e-06, 2.7508431e-06, -3.3284992e-05, -0.00019685866, 5.465961e-06, 2.5712827e-06, -0.0001307662, -0.00019268612, 8.368619e-06, 2.3671205e-06, -0.00022559743, -0.0001862756, 1.111513e-05, 2.1411277e-06, -0.0003166869, -0.00017773996, 1.3676734e-05, 1.896278e-06, -0.00040300505, -0.00016721482, 1.6027298e-05, 1.635709e-06, -0.00048359542, -0.00015485672, 1.814357e-05, 1.3626835e-06, -0.0005575847, -0.00014084089, 2.0005407e-05, 1.0805502e-06, -0.00062419113, -0.00012535887, 2.1595948e-05, 7.927032e-07, -0.0006827326, -0.000108616085, 2.2901751e-05, 5.025426e-07, -0.0007326324, -9.082921e-05, 2.3912902e-05, 2.1343516e-07, -0.0007734245, -7.222342e-05, 2.4623056e-05, -7.132415e-08, -0.00080475706, -5.3029675e-05, 2.502946e-05, -3.4854867e-07, -0.0008263945, -3.3481938e-05, 2.513292e-05, -6.1519495e-07, -0.0008382184, -1.3814398e-05, 2.4937726e-05, -8.6839543e-07, -0.00084022695, 5.7412394e-06, 2.445156e-05, -1.1054885e-06, -0.000832533, 2.4958403e-05, 2.3685325e-05, -1.3240457e-06, -0.0008153609, 4.36182e-05, 2.2652985e-05, -1.5218957e-06, -0.00078904204, 6.151183e-05, 2.1371345e-05, -1.6971446e-06, -0.0007540092, 7.844284e-05, 1.98598e-05, -1.8481938e-06, -0.0007107897, 9.4229166e-05, 1.8140086e-05, -1.973753e-06, -0.0006599982, 0.00010870506, 1.6235963e-05, -2.072849e-06, -0.0006023276, 0.00012172271, 1.4172929e-05, -2.1448332e-06, -0.0005385399, 0.00013315363, 1.197788e-05, -2.189382e-06, -0.0004694564, 0.0001428899, 9.678783e-06, -2.2064958e-06, -0.00039594696, 0.000150845, 7.3043298e-06, -2.1964927e-06, -0.0003189192, 0.00015695447, 4.8835964e-06, -2.16e-06, -0.00023930735, 0.00016117636, 2.4456945e-06, -2.0979417e-06, -0.000158061, 0.00016349126, 1.9438557e-08, -2.0115217e-06, -7.613381e-05, 0.00016390221, -2.3669863e-06, -1.9022065e-06, 5.5276073e-06, 0.00016243423, -4.6863383e-06, -1.7717024e-06, 8.599451e-05, 0.00015913373, -6.91262e-06, -1.6219325e-06, 0.00016436652, 0.00015406757, -9.021357e-06, -1.4550101e-06, 0.0002397816, 0.000147322, -1.09898565e-05, -1.2732113e-06, 0.00031142536, 0.00013900126, -1.2797443e-05, -1.0789458e-06, 0.00037853981, 0.00012922616, -1.4425657e-05, -8.7472654e-07, 0.0004404311, 0.000118132346, -1.585844e-05, -6.631388e-07, 0.0004964765, 0.000105868516, -1.7082273e-05, -4.4680903e-07, 0.0005461306, 9.259446e-05, -1.8086295e-05, -2.2837375e-07, 0.0005889301, 7.847905e-05, -1.8862385e-05, -1.0448686e-08, 0.00062449806, 6.369811e-05, -1.94052e-05, 2.0440125e-07, 0.00065254676, 4.84323e-05, -1.9712208e-05, 4.1369077e-07, 0.0006728795, 3.2864893e-05, -1.9783653e-05, 6.150418e-07, 0.0006853914, 1.7179666e-05, -1.9622514e-05, 8.062092e-07, 0.00069006934, 1.5587267e-06, -1.9234425e-05, 9.851045e-07, 0.00068699016, -1.3819545e-05, -1.8627563e-05, 1.1498179e-06, 0.0006763186, -2.8782508e-05, -1.7812508e-05, 1.2986367e-06, 0.00065830396, -4.316516e-05, -1.6802087e-05, 1.4300626e-06, 0.0006332757, -5.6811925e-05, -1.5611182e-05, 1.5428252e-06, 0.0006016385, -6.957828e-05, -1.4256523e-05, 1.6358925e-06, 0.000563866, -8.1332255e-05, -1.2756469e-05, 1.7084797e-06, 0.00052049453, -9.195575e-05, -1.1130761e-05, 1.7600535e-06, 0.00047211576, -0.00010134568, -9.4002735e-06, 1.7903343e-06, 0.00041936894, -0.00010941489, -7.5867533e-06, 1.7992952e-06, 0.00036293277, -0.000116092924, -5.712553e-06, 1.7871583e-06, 0.00030351683, -0.00012132655, -3.8003616e-06, 1.7543875e-06, 0.00024185305, -0.00012508009, -1.8729359e-06, 1.7016795e-06, 0.00017868665, -0.00012733552, 4.716473e-08, 1.6299514e-06, 0.00011476754, -0.00012809242, 1.9378356e-06, 1.540327e-06, 5.0841467e-05, -0.0001273677, 3.7776758e-06, 1.43412e-06, -1.2358492e-05, -0.00012519505, 5.5462247e-06, 1.3128151e-06, -7.412017e-05, -0.000121624274, 7.224183e-06, 1.1780489e-06, -0.0001337602, -0.00011672055, 8.793616e-06, 1.0315878e-06, -0.00019063136, -0.00011056328, 1.0238141e-05, 8.753053e-07, -0.00024412952, -0.00010324503, 1.154309e-05, 7.1115886e-07, -0.00029369982, -9.487021e-05, 1.269565e-05, 5.4116543e-07, -0.00033884228, -8.555365e-05, 1.3684982e-05, 3.673775e-07, -0.00037911665, -7.541913e-05, 1.4502314e-05, 1.918583e-07, -0.00041414646, -6.459776e-05, 1.5141006e-05, 1.6657985e-08, -0.00044362227, -5.322641e-05, 1.5596595e-05, -1.5621004e-07, -0.00046730423, -4.1445935e-05, 1.5866808e-05, -3.2479178e-07, -0.00048502345, -2.9399558e-05, 1.5951551e-05, -4.872143e-07, -0.000496683, -1.7231143e-05, 1.5852878e-05, -6.417063e-07, -0.00050225767, -5.0835165e-06, 1.5574926e-05, -7.866165e-07, -0.000501793, 6.9031535e-06, 1.5123837e-05, -9.204313e-07, -0.00049540366, 1.8592944e-05, 1.4507653e-05, -1.0417896e-06, -0.00048327097, 2.985567e-05, 1.37361885e-05, -1.1494964e-06, -0.00046563946, 4.0568302e-05, 1.2820891e-05, -1.2425335e-06, -0.00044281324, 5.061626e-05, 1.17746795e-05, -1.3200689e-06, -0.00041515133, 5.989461e-05, 1.0611769e-05, -1.3814628e-06, -0.00038306252, 6.830909e-05, 9.347489e-06, -1.4262722e-06, -0.00034699994, 7.5777054e-05, 7.998085e-06, -1.4542526e-06, -0.00030745493, 8.22282e-05, 6.580511e-06, -1.4653576e-06, -0.0002649508, 8.760522e-05, 5.1122324e-06, -1.4597363e-06, -0.00022003613, 9.186418e-05, 3.6110046e-06, -1.437728e-06, -0.00017327811, 9.4974865e-05, 2.0946684e-06, -1.3998554e-06, -0.00012525555, 9.692086e-05, 5.8094145e-07, -1.3468156e-06, -7.655202e-05, 9.769953e-05, -9.127852e-07, -1.2794687e-06, -2.7749007e-05, 9.732179e-05, -2.3696427e-06, -1.198826e-06, 2.058078e-05, 9.581178e-05, -3.7734703e-06, -1.1060347e-06, 6.7879904e-05, 9.320637e-05, -5.1089905e-06, -1.0023633e-06, 0.000113612405, 8.955446e-05, -6.3619723e-06, -8.8918443e-07, 0.00015726963, 8.491628e-05, -7.5193757e-06, -7.6795754e-07, 0.00019837571, 7.9362464e-05, -8.569485e-06, -6.402103e-07, 0.00023649246, 7.2973075e-05, -9.502019e-06, -5.075201e-07, 0.00027122386, 6.5836495e-05, -1.0308231e-05, -3.7149482e-07, 0.00030221997, 5.8048292e-05, -1.0980981e-05, -2.3375374e-07, 0.0003291801, 4.970997e-05, -1.1514789e-05, -9.590874e-08, 0.0003518556, 4.09277e-05, -1.1905875e-05, 4.045425e-08, 0.0003700517, 3.1811025e-05, -1.2152172e-05, 1.7379317e-07, 0.0003836291, 2.247151e-05, -1.2253321e-05, 3.026269e-07, 0.00039250444, 1.3021434e-05, -1.2210649e-05, 4.2555126e-07, 0.00039665043, 3.5724718e-06, -1.2027122e-05, 5.4125417e-07, 0.00039609513, -5.7655866e-06, -1.1707282e-05, 6.48529e-07, 0.00039092085, -1.488608e-05, -1.1257177e-05, 7.46287e-07, 0.00038126216, -2.3686656e-05, -1.06842535e-05, 8.3356764e-07, 0.00036730347, -3.2070388e-05, -9.997255e-06, 9.095478e-07, 0.00034927618, -3.99468e-05, -9.206096e-06, 9.735488e-07, 0.00032745497, -4.7232814e-05, -8.32173e-06, 1.0250419e-06, 0.00030215413, -5.3853582e-05, -7.3560022e-06, 1.0636519e-06, 0.00027372318, -5.9743223e-05, -6.3214984e-06, 1.0891589e-06, 0.00024254216, -6.484542e-05, -5.231389e-06, 1.1014981e-06, 0.00020901674, -6.911395e-05, -4.0992645e-06, 1.1007583e-06, 0.00017357318, -7.2512994e-05, -2.9389716e-06, 1.0871773e-06, 0.00013665296, -7.501741e-05, -1.7644494e-06, 1.0611384e-06, 9.87074e-05, -7.6612865e-05, -5.895656e-07, 1.0231615e-06, 6.0192346e-05, -7.729579e-05, 5.720419e-07, 9.738964e-07, 2.1562724e-05, -7.707322e-05, 1.70712e-06, 9.141121e-07, -1.6732654e-05, -7.596262e-05, 2.802946e-06, 8.446863e-07, -5.425622e-05, -7.399141e-05, 3.8474677e-06, 7.6659353e-07, -9.058652e-05, -7.119654e-05, 4.82943e-06, 6.808917e-07, -0.00012532285, -6.762388e-05, 5.7384927e-06, 5.887091e-07, -0.0001580895, -6.332756e-05, 6.565335e-06, 4.912297e-07, -0.00018853977, -5.8369184e-05, 7.3017445e-06, 3.8967877e-07, -0.00021635942, -5.2817e-05, 7.940697e-06, 2.8530778e-07, -0.00024126982, -4.6744997e-05, 8.476415e-06, 1.7937968e-07, -0.00026303058, -4.0231964e-05, 8.904414e-06, 7.3153934e-08, -0.00028144172, -3.3360477e-05, 9.221534e-06, -3.2127932e-08, -0.00029634527, -2.6215896e-05, 9.425953e-06, -1.3525641e-07, -0.00030762635, -1.8885325e-05, 9.517186e-06, -2.350675e-07, -0.00031521395, -1.1456575e-05, 9.496067e-06, -3.3045538e-07, -0.0003190809, -4.017131e-06, 9.3647195e-06, -4.2038428e-07, -0.00031924344, 3.3468475e-06, 9.126507e-06, -5.038993e-07, -0.00031576038, 1.0551507e-05, 8.785978e-06, -5.80136e-07, -0.00030873172, 1.7516233e-05, 8.348788e-06, -6.48329e-07, -0.00029829674, 2.4164523e-05, 7.821619e-06, -7.0781925e-07, -0.00028463174, 3.042481e-05, 7.2120833e-06, -7.580597e-07, -0.00026794747, 3.6231206e-05, 6.5286226e-06, -7.9861974e-07, -0.00024848603, 4.152417e-05, 5.7803913e-06, -8.291885e-07, -0.0002265176, 4.625109e-05, 4.9771434e-06, -8.4957605e-07, -0.0002023368, 5.036678e-05, 4.1291064e-06, -8.597141e-07, -0.00017625892, 5.383387e-05, 3.2468565e-06, -8.59654e-07, -0.00014861595, 5.6623125e-05, 2.3411897e-06, -8.4956497e-07, -0.00011975233, 5.8713624e-05, 1.4229928e-06, -8.2972946e-07, -9.002095e-05, 6.0092883e-05, 5.031167e-07, -8.005384e-07, -5.977878e-05, 6.0756858e-05, -4.0774938e-07, -7.624847e-07, -2.9382736e-05, 6.0709834e-05, -1.2991989e-06, -7.161559e-07, 8.14462e-07, 5.9964248e-05, -2.1612236e-06, -6.622257e-07, 3.0468289e-05, 5.8540416e-05, -2.9843227e-06, -6.0144475e-07, 5.9246275e-05, 5.6466146e-05, -3.7596046e-06, -5.346306e-07, 8.6831635e-05, 5.377632e-05, -4.4788794e-06, -4.6265728e-07, 0.000112926675, 5.0512335e-05, -5.1347433e-06, -3.86444e-07, 0.00013725593, 4.6721547e-05, -5.7206485e-06, -3.0694392e-07, 0.00015956897, 4.2456617e-05, -6.230967e-06, -2.2513252e-07, 0.00017964284, 3.777479e-05, -6.6610396e-06, -1.4199584e-07, 0.00019728423, 3.2737193e-05, -7.0072147e-06, -5.8518935e-08, 0.0002123312, 2.7408027e-05, -7.2668718e-06, 2.4325521e-08, 0.00022465452, 2.1853803e-05, -7.438435e-06, 1.0558829e-07, 0.00023415861, 1.6142507e-05, -7.5213766e-06, 1.8435419e-07, 0.00024078209, 1.0342813e-05, -7.516201e-06, 2.597521e-07, 0.0002444979, 4.523257e-06, -7.4244263e-06, 3.3096438e-07, 0.0002453131, -1.2485418e-06, -7.2485464e-06, 3.9723534e-07, 0.00024326815, -6.9066514e-06, -6.991987e-06, 4.5787905e-07, 0.00023843585, -1.2387563e-05, -6.6590515e-06, 5.1228614e-07, 0.00023092006, -1.7630884e-05, -6.2548543e-06, 5.599294e-07, 0.0002208539, -2.2579985e-05, -5.7852503e-06, 6.0036876e-07, 0.00020839775, -2.718259e-05, -5.256753e-06, 6.3325484e-07, 0.0001937369, -3.139131e-05, -4.676449e-06, 6.583313e-07, 0.00017707904, -3.516412e-05, -4.051906e-06, 6.754366e-07, 0.00015865147, -3.846473e-05, -3.3910783e-06, 6.84504e-07, 0.00013869806, -4.1262923e-05, -2.702206e-06, 6.8556096e-07, 0.00011747629, -4.3534823e-05, -1.9937172e-06, 6.78727e-07, 9.5253905e-05, -4.526303e-05, -1.274126e-06, 6.642111e-07, 7.2305746e-05, -4.6436733e-05, -5.5193306e-07, 6.423075e-07, 4.891038e-05, -4.705172e-05, 1.6447315e-07, 6.133911e-07, 2.5346864e-05, -4.7110312e-05, 8.6691074e-07, 5.779116e-07, 1.8914722e-06, -4.662124e-05, 1.5474963e-06, 5.363872e-07, -2.1185442e-05, -4.559942e-05, 2.1987307e-06, 4.893973e-07, -4.3622476e-05, -4.4065688e-05, 2.81358e-06, 4.375749e-07, -6.517005e-05, -4.204645e-05, 3.3855483e-06, 3.815984e-07, -8.55931e-05, -3.9573297e-05, 3.9087445e-06, 3.2218284e-07, -0.00010467357, -3.668254e-05, 4.37794e-06, 2.6007118e-07, -0.00012221262, -3.341471e-05, 4.788619e-06, 1.9602507e-07, -0.00013803263, -2.9814035e-05, 5.137018e-06, 1.3081595e-07, -0.00015197888, -2.5927835e-05, 5.420156e-06, 6.521575e-08, -0.000163921, -2.1805956e-05, 5.6358576e-06, -1.1952672e-11, -0.000173754, -1.7500131e-05, 5.7827638e-06, -6.4120634e-08, -0.00018139913, -1.3063353e-05, 5.860334e-06, -1.263892e-07, -0.0001868043, -8.549245e-06, 5.8688393e-06, -1.8612985e-07, -0.00018994427, -4.011421e-06, 5.8093447e-06, -2.4269556e-07, -0.00019082046, 4.971275e-07, 5.683684e-06, -2.9548684e-07, -0.00018946052, 4.924638e-06, 5.494426e-06, -3.4395785e-07, -0.00018591754, 9.221154e-06, 5.2448327e-06, -3.8762184e-07, -0.00018026902, 1.3339076e-05, 4.9388077e-06, -4.2605583e-07, -0.0001726156, 1.7233668e-05, 4.580844e-06, -4.589044e-07, -0.00016307941, 2.0863534e-05, 4.1759586e-06, -4.8588265e-07, -0.00015180242, 2.4191033e-05, 3.7296281e-06, -5.0677835e-07, -0.00013894434, 2.7182663e-05, 3.2477167e-06, -5.214532e-07, -0.00012468056, 2.9809366e-05, 2.7364015e-06, -5.2984313e-07, -0.00010919985, 3.2046803e-05, 2.202096e-06, -5.319579e-07, -9.27019e-05, 3.3875545e-05, 1.651373e-06, -5.278795e-07, -7.5394855e-05, 3.5281228e-05, 1.090884e-06, -5.177603e-07, -5.7492776e-05, 3.625462e-05, 5.272819e-07, -5.018201e-07, -3.921303e-05, 3.679166e-05, -3.285569e-08, -4.803421e-07, -2.0773752e-05, 3.6893394e-05, -5.83102e-07, -4.5366892e-07, -2.3912733e-06, 3.6565907e-05, -1.1172526e-06, -4.221975e-07, 1.5722333e-05, 3.5820143e-05, -1.6293935e-06, -3.8637359e-07, 3.336164e-05, 3.4671713e-05, -2.113965e-06, -3.466858e-07, 5.033014e-05, 3.3140623e-05, -2.5658196e-06, -3.0365925e-07, 6.644237e-05, 3.1250976e-05, -2.9802754e-06, -2.5784885e-07, 8.152586e-05, 2.9030636e-05, -3.3531614e-06, -2.0983232e-07, 9.542295e-05, 2.6510814e-05, -3.6808583e-06, -1.6020327e-07, 0.00010799231, 2.3725677e-05, -3.960331e-06, -1.0956389e-07, 0.00011911037, 2.0711894e-05, -4.189153e-06, -5.8517998e-08, 0.0001286724, 1.750816e-05, -4.365525e-06, -7.663899e-09, 0.00013659344, 1.41547325e-05, -4.488286e-06, 4.2412374e-08, 0.00014280893, 1.0692924e-05, -4.556914e-06, 9.114367e-08, 0.00014727515, 7.1646145e-06, -4.5715233e-06, 1.3798794e-07, 0.00014996933, 3.6117533e-06, -4.5328516e-06, 1.8243412e-07, 0.00015088962, 7.587294e-08, -4.4422413e-06, 2.2400754e-07, 0.00015005471, -3.4023838e-06, -4.301613e-06, 2.622747e-07, 0.0001475033, -6.7837195e-06, -4.1134344e-06, 2.968478e-07, 0.00014329332, -1.0030616e-05, -3.880684e-06, 3.2738822e-07, 0.00013750092, -1.3107738e-05, -3.6068036e-06, 3.536098e-07, 0.00013021928, -1.5982303e-05, -3.2956561e-06, 3.752812e-07, 0.00012155731, -1.8624423e-05, -2.9514704e-06, 3.9222766e-07, 0.00011163802, -2.1007401e-05, -2.5787865e-06, 4.043321e-07, 0.00010059696, -2.3107985e-05, -2.182399e-06, 4.1153544e-07, 8.8580375e-05, -2.4906572e-05, -1.7672962e-06, 4.138364e-07, 7.574336e-05, -2.6387395e-05, -1.3386002e-06, 4.1129053e-07, 6.2247935e-05, -2.7538621e-05, -9.0150434e-07, 4.0400852e-07, 4.826102e-05, -2.8352426e-05, -4.6121215e-07, 3.9215408e-07, 3.395243e-05, -2.8825028e-05, -2.2877371e-08, 3.759412e-07, 1.9492882e-05, -2.8956656e-05, 4.0845538e-07, 3.5563068e-07, 5.0519816e-06, -2.8751478e-05, 8.279069e-07, 3.315265e-07, -9.203712e-06, -2.8217493e-05, 1.2308172e-06, 3.0397143e-07, -2.3112565e-05, -2.7366372e-05, 1.6127958e-06, 2.7334247e-07, -3.6519654e-05, -2.6213258e-05, 1.9697682e-06, 2.4004595e-07, -4.9278453e-05, -2.4776538e-05, 2.298017e-06, 2.045123e-07, -6.125238e-05, -2.3077575e-05, 2.5942204e-06, 1.6719062e-07, -7.2316216e-05, -2.1140404e-05, 2.8554823e-06, 1.2854323e-07, -8.2357365e-05, -1.8991419e-05, 3.0793606e-06, 8.904007e-08, -9.127695e-05, -1.6659023e-05, 3.2638857e-06, 4.9153147e-08, -9.899071e-05, -1.4173269e-05, 3.4075777e-06, 9.350997e-09, -0.00010542977, -1.1565476e-05, 3.509453e-06, -2.9906634e-08, -0.000110541114, -8.8678535e-06, 3.5690296e-06, -6.8173996e-08, -0.000114288, -6.113115e-06, 3.5863227e-06, -1.05024256e-07, -0.00011665008, -3.3340827e-06, 3.561837e-06, -1.4005413e-07, -0.00011762337, -5.6331345e-07, 3.4965524e-06, -1.7288812e-07, -0.000117220006, 2.1672777e-06, 3.3919043e-06, -2.0318245e-07, -0.00011546787, 4.826775e-06, 3.2497605e-06, -2.306285e-07, -0.00011240995, 7.3856017e-06, 3.0723913e-06, -2.5495575e-07, -0.00010810364, 9.815843e-06, 2.8624365e-06, -2.7593435e-07, -0.00010261982, 1.2091539e-05, 2.6228697e-06, -2.9337704e-07, -9.604178e-05, 1.4188953e-05, 2.3569569e-06, -3.071406e-07, -8.8464105e-05, 1.608681e-05, 2.0682148e-06, -3.1712682e-07, -7.9991325e-05, 1.7766497e-05, 1.7603655e-06, -3.2328285e-07, -7.07366e-05, 1.9212242e-05, 1.4372904e-06, -3.256011e-07, -6.0820214e-05, 2.0411244e-05, 1.1029816e-06, -3.2411845e-07, -5.0368115e-05, 2.1353771e-05, 7.6149513e-07, -3.1891526e-07, -3.951032e-05, 2.203322e-05, 4.1690186e-07, -3.1011356e-07, -2.8379354e-05, 2.244615e-05, 7.3240784e-08, -2.97875e-07, -1.7108689e-05, 2.2592254e-05, -2.6552746e-07, -2.8239836e-07, -5.8311625e-06, 2.2474325e-05, -5.955651e-07, -2.6391652e-07, 5.322533e-06, 2.209816e-05, -9.131995e-07, -2.426933e-07, 1.6225336e-05, 2.1472451e-05, -1.2149629e-06, -2.1901977e-07, 2.6755224e-05, 2.0608632e-05, -1.4976296e-06, -1.9321064e-07, 3.6796537e-05, 1.95207e-05, -1.7582483e-06, -1.6559994e-07, 4.6241214e-05, 1.8225011e-05, -1.9941729e-06, -1.3653707e-07, 5.4989916e-05, 1.6740056e-05, -2.2030865e-06, -1.0638233e-07, 6.295303e-05, 1.5086201e-05, -2.3830241e-06, -7.550269e-08, 7.0051545e-05, 1.32854275e-05, -2.532389e-06, -4.4267367e-08, 7.621777e-05, 1.1361051e-05, -2.649965e-06, -1.3043507e-08, 8.139596e-05, 9.337426e-06, -2.7349233e-06, 1.7807992e-08, 8.554275e-05, 7.2396447e-06, -2.786828e-06, 4.7936574e-08, 8.862743e-05, 5.0932417e-06, -2.8056313e-06, 7.7005915e-08, 9.063209e-05, 2.9238838e-06, -2.7916708e-06, 1.04697556e-07, 9.1551665e-05, 7.5707374e-07, -2.7456565e-06, 1.3071431e-07, 9.1393704e-05, -1.3821424e-06, -2.6686582e-06, 1.5478335e-07, 9.017812e-05, -3.4694579e-06, -2.5620861e-06, 1.7665892e-07, 8.793673e-05, -5.481574e-06, -2.4276687e-06, 1.9612479e-07, 8.47127e-05, -7.396453e-06, -2.2674285e-06, 2.129962e-07, 8.055987e-05, -9.193553e-06, -2.0836526e-06, 2.271215e-07, 7.5541895e-05, -1.0854037e-05, -1.8788618e-06, 2.3838341e-07, 6.97314e-05, -1.2360969e-05, -1.6557786e-06, 2.4669964e-07, 6.320899e-05, -1.3699472e-05, -1.4172914e-06, 2.5202348e-07, 5.6062112e-05, -1.4856868e-05, -1.1664183e-06, 2.5434352e-07, 4.8384034e-05, -1.5822789e-05, -9.0627026e-07, 2.5368337e-07, 4.0272582e-05, -1.6589256e-05, -6.400135e-07, 2.501007e-07, 3.1828968e-05, -1.7150733e-05, -3.7083197e-07, 2.4368606e-07, 2.3156555e-05, -1.7504153e-05, -1.01890066e-07, 2.3456117e-07, 1.435963e-05, -1.7648905e-05, 1.6370362e-07, 2.2287718e-07, 5.5421697e-06, -1.7586804e-05, 4.229313e-07, 2.0881225e-07, -3.1933469e-06, -1.7322034e-05, 6.728994e-07, 1.9256915e-07, -1.1747107e-05, -1.686105e-05, 9.108701e-07, 1.743724e-07, -2.0023072e-05, -1.621247e-05, 1.1342902e-06, 1.5446543e-07, -2.7930024e-05, -1.5386946e-05, 1.3408177e-06, 1.3310733e-07, -3.5382545e-05, -1.4396995e-05, 1.5283455e-06, 1.1056968e-07, -4.2301916e-05, -1.32568275e-05, 1.6950215e-06, 8.7133124e-08, -4.861689e-05, -1.1982159e-05, 1.8392662e-06, 6.3084016e-08, -5.4264423e-05, -1.0589995e-05, 1.9597862e-06, 3.8711e-08, -5.9190246e-05, -9.0984195e-06, 2.0555842e-06, 1.430163e-08, -6.334936e-05, -7.5263633e-06, 2.1259661e-06, -9.860944e-09, -6.670639e-05, -5.893373e-06, 2.170543e-06, -3.350118e-08, -6.923584e-05, -4.219372e-06, 2.189232e-06, -5.6354196e-08, -7.092221e-05, -2.5244262e-06, 2.1822507e-06, -7.816867e-08, -7.176004e-05, -8.285087e-07, 2.1501103e-06, -9.8709506e-08, -7.175378e-05, 8.4873153e-07, 2.093605e-06, -1.1776031e-07, -7.091756e-05, 2.48819e-06, 2.0137973e-06, -1.3512555e-07, -6.92749e-05, 4.071519e-06, 1.9120018e-06, -1.5063247e-07, -6.685826e-05, 5.5813275e-06, 1.7897659e-06, -1.6413277e-07, -6.370851e-05, 7.0013675e-06, 1.648847e-06, -1.7550381e-07, -5.987432e-05, 8.316701e-06, 1.4911902e-06, -1.8464969e-07, -5.541149e-05, 9.513851e-06, 1.318901e-06, -1.9150185e-07, -5.038214e-05, 1.0580937e-05, 1.1342196e-06, -1.9601949e-07, -4.485392e-05, 1.150778e-05, 9.3949166e-07, -1.9818941e-07, -3.8899136e-05, 1.22859965e-05, 7.371402e-07, -1.9802593e-07, -3.2593794e-05, 1.2909061e-05, 5.296358e-07, -1.9557007e-07, -2.6016718e-05, 1.3372358e-05, 3.1946735e-07, -1.9088873e-07, -1.9248537e-05, 1.3673193e-05, 1.09112754e-07, -1.8407341e-07, -1.2370756e-05, 1.3810802e-05, -9.898927e-08, -1.7523885e-07, -5.4647835e-06, 1.3786319e-05, -3.0246696e-07, -1.645212e-07, 1.3890079e-06, 1.3602737e-05, -4.9904185e-07, -1.5207614e-07, 8.1121925e-06, 1.3264842e-05, -6.8655345e-07, -1.3807673e-07, 1.4629167e-05, 1.2779124e-05, -8.6298246e-07, -1.2271113e-07, 2.086798e-05, 1.2153676e-05, -1.0264716e-06, -1.0618019e-07, 2.67611e-05, 1.1398073e-05, -1.1753446e-06, -8.869485e-08, 3.2246127e-05, 1.05232375e-05, -1.3081221e-06, -7.047359e-08, 3.726643e-05, 9.541287e-06, -1.4235364e-06, -5.1739743e-08, 4.1771702e-05, 8.4653775e-06, -1.5205416e-06, -3.2718837e-08, 4.5718432e-05, 7.309533e-06, -1.5983226e-06, -1.36359475e-08, 4.907031e-05, 6.0884668e-06, -1.6563004e-06, 5.286898e-09, 5.1798514e-05, 4.8174015e-06, -1.6941349e-06, 2.3833246e-08, 5.388192e-05, 3.511883e-06, -1.711725e-06, 4.1794628e-08, 5.530722e-05, 2.1875971e-06, -1.7092055e-06, 5.8972827e-08, 5.606895e-05, 8.601836e-07, -1.6869421e-06, 7.518202e-08, 5.616941e-05, -4.5494357e-07, -1.6455224e-06, 9.0250715e-08, 5.561852e-05, -1.7427701e-06, -1.5857463e-06, 1.04023485e-07, 5.4433567e-05, -2.9888492e-06, -1.5086126e-06, 1.16362514e-07, 5.2638887e-05, -4.179459e-06, -1.4153046e-06, 1.2714888e-07, 5.026547e-05, -5.3017493e-06, -1.3071726e-06, 1.3628365e-07, 4.735048e-05, -6.343876e-06, -1.1857163e-06, 1.4368864e-07, 4.393673e-05, -7.29512e-06, -1.0525642e-06, 1.49307e-07, 4.0072082e-05, -8.145996e-06, -9.094535e-07, 1.5310354e-07, 3.580882e-05, -8.888336e-06, -7.582069e-07, 1.5506474e-07, 3.1202966e-05, -9.515367e-06, -6.0071125e-07, 1.5519853e-07, 2.6313564e-05, -1.0021764e-05, -4.3889403e-07, 1.535339e-07, 2.1201959e-05, -1.0403686e-05, -2.7470048e-07, 1.5012013e-07, 1.5931031e-05, -1.0658799e-05, -1.100708e-07, 1.4502596e-07, 1.0564455e-05, -1.0786274e-05, 5.3082175e-08, 1.3833844e-07, 5.1659445e-06, -1.07867745e-05, 2.1289476e-07, 1.3016155e-07, -2.0148215e-07, -1.0662422e-05, 3.675731e-07, 1.2061484e-07, -5.4762245e-06, -1.0416747e-05, 5.1541275e-07, 1.0983168e-07, -1.0598786e-05, -1.0054626e-05, 6.548171e-07, 9.795754e-08, -1.5512429e-05, -9.5822015e-06, 7.843136e-07, 8.514806e-08, -2.0163783e-05, -9.00679e-06, 9.025693e-07, 7.156713e-08, -2.450341e-05, -8.336776e-06, 1.0084035e-06, 5.7384813e-08, -2.8486307e-05, -7.5815014e-06, 1.1007993e-06, 4.2775305e-08, -3.2072356e-05, -6.7511364e-06, 1.1789118e-06, 2.7914819e-08, -3.5226698e-05, -5.8565506e-06, 1.2420762e-06, 1.29795295e-08, -3.7920065e-05, -4.9091745e-06, 1.2898115e-06, -1.8564684e-09, -4.012901e-05, -3.9208594e-06, 1.3218233e-06, -1.6423142e-08, -4.1836083e-05, -2.9037305e-06, 1.3380044e-06, -3.0556418e-08, -4.302994e-05, -1.8700448e-06, 1.3384324e-06, -4.4099988e-08, -4.370537e-05, -8.320446e-07, 1.3233658e-06, -5.6906977e-08, -4.386325e-05, 1.9818224e-07, 1.2932386e-06, -6.8841494e-08, -4.3510423e-05, 1.2088404e-06, 1.2486513e-06, -7.978004e-08, -4.265954e-05, 2.1885587e-06, 1.1903622e-06, -8.961266e-08, -4.1328803e-05, 3.1265147e-06, 1.1192752e-06, -9.82441e-08, -3.954166e-05, 4.01255e-06, 1.0364272e-06, -1.0559456e-07, -3.7326456e-05, 4.837278e-06, 9.42974e-07, -1.1160041e-07, -3.471601e-05, 5.5921782e-06, 8.4017483e-07, -1.1621466e-07, -3.1747168e-05, 6.269682e-06, 7.293758e-07, -1.1940719e-07, -2.8460314e-05, 6.863243e-06, 6.1199336e-07, -1.2116487e-07, -2.4898829e-05, 7.367396e-06, 4.8949624e-07, -1.2149137e-07, -2.1108548e-05, 7.777802e-06, 3.633879e-07, -1.2040688e-07, -1.713719e-05, 8.0912805e-06, 2.3518831e-07, -1.17947565e-07, -1.3033769e-05, 8.305825e-06, 1.0641632e-07, -1.14164905e-07, -8.848008e-06, 8.42061e-06, -2.1428088e-08, -1.0912485e-07, -4.6297487e-06, 8.435976e-06, -1.4688077e-07, -1.02906775e-07, -4.283758e-07, 8.353412e-06, -2.6852976e-07, -9.5602374e-08, 3.7077489e-06, 8.1755115e-06, -3.8503077e-07, -8.731437e-08, 7.731828e-06, 7.905931e-06, -4.9512164e-07, -7.815517e-08, 1.1599147e-05, 7.5493263e-06, -5.9763545e-07, -6.824535e-08, 1.5267551e-05, 7.1112827e-06, -6.9151264e-07, -5.7712192e-08, 1.8697896e-05, 6.5982344e-06, -7.758113e-07, -4.668803e-08, 2.1854452e-05, 6.0173766e-06, -8.497161e-07, -3.5308684e-08, 2.4705249e-05, 5.3765684e-06, -9.125458e-07, -2.3711806e-08, 2.7222399e-05, 4.6842315e-06, -9.637586e-07, -1.2035253e-08, 2.938234e-05, 3.949244e-06, -1.0029563e-06, -4.1550688e-10, 3.1166037e-05, 3.1808268e-06, -1.0298866e-06, 1.10139e-08, 3.255914e-05, 2.3884359e-06, -1.0444431e-06, 2.2123873e-08, 3.3552045e-05, 1.5816453e-06, -1.0466648e-06, 3.2791178e-08, 3.4139954e-05, 7.7003534e-07, -1.0367326e-06, 4.2899764e-08, 3.432283e-05, -3.69178e-08, -1.0149648e-06, 5.2341996e-08, 3.410533e-05, -8.2995075e-07, -9.818118e-07, 6.1019755e-08, 3.349667e-05, -1.6001162e-06, -9.378482e-07, 6.88454e-08, 3.251043e-05, -2.3388816e-06, -8.8376385e-07, 7.574265e-08, 3.1164345e-05, -3.03822e-06, -8.2035433e-07, 8.1647215e-08, 2.948001e-05, -3.6906963e-06, -7.485099e-07, 8.650739e-08, 2.7482578e-05, -4.2895413e-06, -6.692034e-07, 9.028442e-08, 2.5200407e-05, -4.82872e-06, -5.83478e-07, 9.295275e-08, 2.2664673e-05, -5.3029903e-06, -4.9243346e-07, 9.450006e-08, 1.9908968e-05, -5.707948e-06, -3.972128e-07, 9.492723e-08, 1.696887e-05, -6.0400644e-06, -2.9898823e-07, 9.424809e-08, 1.3881489e-05, -6.2967147e-06, -1.989471e-07, 9.248904e-08, 1.0685027e-05, -6.4761903e-06, -9.827793e-08, 8.968854e-08, 7.4183044e-06, -6.5777053e-06, 1.8434313e-09, 8.589646e-08, 4.120308e-06, -6.6013895e-06, 1.0026714e-07, 8.117331e-08, 8.2973276e-07, -6.54827e-06, 1.9588225e-07, 7.558938e-08, -2.4154588e-06, -6.4202472e-06, 2.8762895e-07, 6.9223724e-08, -5.5784653e-06, -6.220056e-06, 3.7450994e-07, 6.216313e-08, -8.624052e-06, -5.951222e-06, 4.5560094e-07, 5.4500983e-08, -1.1518933e-05, -5.618005e-06, 5.3006016e-07, 4.6336062e-08, -1.4232124e-05, -5.225339e-06, 5.971367e-07, 3.777131e-08, -1.6735263e-05, -4.7787644e-06, 6.5617763e-07, 2.8912583e-08, -1.900289e-05, -4.2843517e-06, 7.0663407e-07, 1.9867352e-08, -2.1012702e-05, -3.7486245e-06, 7.4806553e-07, 1.0743461e-08, -2.2745751e-05, -3.178475e-06, 7.801436e-07, 1.6478545e-09, -2.4186611e-05, -2.5810787e-06, 8.026534e-07, -7.314643e-09, -2.5323492e-05, -1.9638057e-06, 8.1549456e-07, -1.6042502e-08, -2.6148327e-05, -1.334134e-06, 8.186803e-07, -2.4438608e-08, -2.6656788e-05, -6.99559e-07, 8.1233526e-07, -3.2411315e-08, -2.6848285e-05, -6.750777e-08, 7.966925e-07, -3.987541e-08, -2.672591e-05, 5.5474624e-07, 7.7208864e-07, -4.6752994e-08, -2.629633e-05, 1.1601646e-06, 7.3895853e-07, -5.297427e-08, -2.5569658e-05, 1.7420219e-06, 6.9782834e-07, -5.8478193e-08, -2.4559278e-05, 2.2939776e-06, 6.493081e-07, -6.321305e-08, -2.3281635e-05, 2.8101433e-06, 5.940831e-07, -6.713691e-08, -2.1755988e-05, 3.2851442e-06, 5.3290483e-07, -7.021791e-08, -2.0004149e-05, 3.7141713e-06, 4.665811e-07, -7.243448e-08, -1.8050176e-05, 4.093028e-06, 3.9596574e-07, -7.377544e-08, -1.5920072e-05, 4.4181697e-06, 3.21948e-07, -7.42399e-08, -1.3641439e-05, 4.686732e-06, 2.454416e-07, -7.3837164e-08, -1.1243135e-05, 4.8965535e-06, 1.6737378e-07, -7.2586396e-08, -8.754923e-06, 5.046189e-06, 8.8674355e-08, -7.0516265e-08, -6.2071076e-06, 5.134914e-06, 1.0264847e-08, -6.766444e-08, -3.630174e-06, 5.162721e-06, -6.6951976e-08, -6.407701e-08, -1.0544359e-06, 5.1303095e-06, -1.4210227e-07, -5.980781e-08, 1.4903147e-06, 5.0390613e-06, -2.1435072e-07, -5.4917674e-08, 3.9751435e-06, 4.8910183e-06, -2.829096e-07, -4.947358e-08, 6.3722937e-06, 4.6888445e-06, -3.4704712e-07, -4.354783e-08, 8.655489e-06, 4.435787e-06, -4.060948e-07, -3.721706e-08, 1.08002105e-05, 4.1356266e-06, -4.594544e-07, -3.056134e-08, 1.2783956e-05, 3.792626e-06, -5.0660344e-07, -2.3663135e-08, 1.4586458e-05, 3.411473e-06, -5.471001e-07, -1.660636e-08, 1.6189892e-05, 2.9972182e-06, -5.8058697e-07, -9.475348e-09, 1.757903e-05, 2.5552106e-06, -6.067938e-07, -2.3538813e-09, 1.8741386e-05, 2.091031e-06, -6.2553903e-07, 4.675767e-09, 1.9667305e-05, 1.6104239e-06, -6.3673053e-07, 1.1533766e-08, 2.0350028e-05, 1.1192269e-06, -6.403653e-07, 1.8143606e-08, 2.0785727e-05, 6.233033e-07, -6.365276e-07, 2.4432934e-08, 2.0973497e-05, 1.2847242e-07, -6.2538703e-07, 3.0334313e-08, 2.0915319e-05, -3.5955634e-07, -6.071947e-07, 3.5785927e-08, 2.0615984e-05, -8.3524793e-07, -5.8227926e-07, 4.0732203e-08, 2.0082998e-05, -1.2933027e-06, -5.510416e-07, 4.512434e-08, 1.9326444e-05, -1.7287141e-06, -5.139491e-07, 4.8920786e-08, 1.8358827e-05, -2.136821e-06, -4.7152912e-07, 5.208755e-08, 1.719488e-05, -2.513357e-06, -4.2436182e-07, 5.459853e-08, 1.5851365e-05, -2.854492e-06, -3.730726e-07, 5.6435628e-08, 1.4346844e-05, -3.1568707e-06, -3.1832414e-07, 5.7588863e-08, 1.2701429e-05, -3.417641e-06, -2.6080804e-07, 5.805633e-08, 1.0936526e-05, -3.6344818e-06, -2.0123633e-07, 5.784409e-08, 9.074568e-06, -3.8056182e-06, -1.40333e-07, 5.6965984e-08, 7.138734e-06, -3.9298347e-06, -7.882523e-08, 5.544332e-08, 5.152669e-06, -4.0064797e-06, -1.7435102e-08, 5.33045e-08, 3.1402064e-06, -4.0354616e-06, 4.312879e-08, 5.0584603e-08, 1.1250844e-06, -4.0172436e-06, 1.02179264e-07, 4.7324832e-08, -8.693256e-07, -3.9528263e-06, 1.5905817e-07, 4.3571955e-08, -2.8202828e-06, -3.8437292e-06, 2.131435e-07, 3.937766e-08, -4.70593e-06, -3.6919637e-06, 2.6385598e-07, 3.4797885e-08, -6.5055324e-06, -3.5000005e-06, 3.1066514e-07, 2.9892096e-08, -8.199699e-06, -3.2707346e-06, 3.530945e-07, 2.4722523e-08, -9.770581e-06, -3.0074448e-06, 3.9072623e-07, 1.935342e-08, -1.120206e-05, -2.713748e-06, 4.2320514e-07, 1.3850275e-08, -1.2479897e-05, -2.3935534e-06, 4.5024154e-07, 8.279025e-09, -1.3591873e-05, -2.0510108e-06, 4.7161362e-07, 2.705293e-09, -1.4527891e-05, -1.6904595e-06, 4.8716885e-07, -2.8063643e-09, -1.5280062e-05, -1.3163748e-06, 4.9682455e-07, -8.193193e-09, -1.5842756e-05, -9.3331323e-07, 5.005677e-07, -1.3394932e-08, -1.6212629e-05, -5.4585934e-07, 4.984541e-07, -1.8354473e-08, -1.6388629e-05, -1.585717e-07, 4.906061e-07, -2.3018469e-08, -1.6371963e-05, 2.2406947e-07, 4.772107e-07, -2.7337883e-08, -1.6166048e-05, 5.9771264e-07, 4.5851576e-07, -3.1268492e-08, -1.5776437e-05, 9.581833e-07, 4.3482646e-07, -3.4771308e-08, -1.5210711e-05, 1.3015293e-06, 4.0650062e-07, -3.781295e-08, -1.447837e-05, 1.624063e-06, 3.7394372e-07, -4.036594e-08, -1.3590677e-05, 1.9223992e-06, 3.376035e-07, -4.2408903e-08, -1.2560508e-05, 2.1934895e-06, 2.9796394e-07, -4.392674e-08, -1.1402173e-05, 2.434652e-06, 2.5553908e-07, -4.4910674e-08, -1.0131225e-05, 2.6435964e-06, 2.1086669e-07, -4.5358256e-08, -8.76426e-06, 2.818443e-06, 1.6450147e-07, -4.527329e-08, -7.31871e-06, 2.9577386e-06, 1.1700846e-07, -4.4665676e-08, -5.8126207e-06, 3.060466e-06, 6.895629e-08, -4.35512e-08, -4.26444e-06, 3.1260481e-06, 2.0910543e-08, -4.195125e-08, -2.692793e-06, 3.1543477e-06, -2.6572744e-08, -3.9892477e-08, -1.1162645e-06, 3.1456611e-06, -7.295335e-08, -3.7406398e-08, 4.4681502e-07, 3.100708e-06, -1.17712865e-07, -3.452894e-08, 1.9785773e-06, 3.0206158e-06, -1.6036032e-07, -3.1299972e-08, 3.4618163e-06, 2.9068997e-06, -2.0043741e-07, -2.7762754e-08, 4.8801753e-06, 2.7614387e-06, -2.3752328e-07, -2.3963391e-08, 6.2183217e-06, 2.586448e-06, -2.712387e-07, -1.9950253e-08, 7.4621094e-06, 2.3844475e-06, -3.0124983e-07, -1.5773377e-08, 8.59872e-06, 2.1582275e-06, -3.2727132e-07, -1.148385e-08, 9.616792e-06, 1.9108118e-06, -3.4906873e-07, -7.133216e-09, 1.0506524e-05, 1.645419e-06, -3.6646045e-07, -2.772857e-09, 1.12597645e-05, 1.3654222e-06, -3.7931895e-07, 1.5465892e-09, 1.1870081e-05, 1.0743067e-06, -3.8757128e-07, 5.7758074e-09, 1.23328e-05, 7.756284e-07, -3.91199e-07, 9.867353e-09, 1.2645036e-05, 4.72971e-07, -3.9023757e-07, 1.3776168e-08, 1.2805693e-05, 1.6990451e-07, -3.8477492e-07, 1.7460064e-08, 1.2815448e-05, -1.3005625e-07, -3.7494965e-07, 2.0880165e-08, 1.2676715e-05, -4.234912e-07, -3.6094852e-07, 2.4001295e-08, 1.2393585e-05, -7.07113e-07, -3.4300348e-07, 2.6792332e-08, 1.19717515e-05, -9.77803e-07, -3.213883e-07, 2.9226493e-08, 1.1418419e-05, -1.2326444e-06, -2.9641464e-07, 3.1281576e-08, 1.0742192e-05, -1.4689527e-06, -2.6842778e-07, 3.294014e-08, 9.952956e-06, -1.6843028e-06, -2.3780213e-07, 3.418962e-08, 9.061738e-06, -1.8765529e-06, -2.0493634e-07, 3.5022403e-08, 8.0805585e-06, -2.0438645e-06, -1.7024837e-07, 3.543582e-08, 7.022283e-06, -2.1847181e-06, -1.3417024e-07, 3.5432116e-08, 5.90045e-06, -2.2979264e-06, -9.714284e-08, 3.5018306e-08, 4.7291087e-06, -2.382642e-06, -5.961066e-08, 3.420605e-08, 3.522645e-06, -2.4383608e-06, -2.201661e-08, 3.3011418e-08, 2.2956121e-06, -2.4649235e-06, 1.5203117e-08, 3.145464e-08, 1.0625567e-06, -2.4625108e-06, 5.1623957e-08, 2.95598e-08, -1.6214814e-07, -2.4316355e-06, 8.68377e-08, 2.7354488e-08, -1.3644666e-06, -2.3731318e-06, 1.2045693e-07, 2.486943e-08, -2.5308568e-06, -2.2881388e-06, 1.5211921e-07, 2.2138071e-08, -3.6484198e-06, -2.1780843e-06, 1.8149078e-07, 1.9196154e-08, -4.7050376e-06, -2.0446614e-06, 2.0827e-07, 1.6081255e-08, -5.6894996e-06, -1.8898058e-06, 2.3219027e-07, 1.2832329e-08, -6.59162e-06, -1.7156688e-06, 2.530226e-07, 9.489224e-09, -7.402335e-06, -1.5245887e-06, 2.7057752e-07, 6.0922143e-09, -8.113791e-06, -1.319061e-06, 2.847067e-07, 2.6815246e-09, -8.719416e-06, -1.1017064e-06, 2.953039e-07, -7.031364e-10, -9.21397e-06, -8.75239e-07, 3.0230558e-07, -4.023026e-09, -9.593588e-06, -6.4243255e-07, 3.0569092e-07, -7.240799e-09, -9.855804e-06, -4.0608802e-07, 3.0548125e-07, -1.0320919e-08, -9.999545e-06, -1.6900032e-07, 3.0173916e-07, -1.3230036e-08, -1.0025133e-05, 6.6073824e-08, 2.945671e-07, -1.5937339e-08, -9.934248e-06, 2.964471e-07, 2.841055e-07, -1.8414866e-08, -9.729894e-06, 5.195316e-07, 2.7053053e-07, -2.0637788e-08, -9.416336e-06, 7.328672e-07, 2.5405143e-07, -2.2584635e-08, -8.999032e-06, 9.3414764e-07, 2.3490755e-07, -2.423749e-08, -8.484549e-06, 1.121245e-06, 2.1336508e-07, -2.5582146e-08, -7.88047e-06, 1.2922309e-06, 1.8971357e-07, -2.6608195e-08, -7.195287e-06, 1.445396e-06, 1.6426205e-07, -2.7309092e-08, -6.4382893e-06, 1.5792658e-06, 1.3733528e-07, -2.7682168e-08, -5.6194417e-06, 1.6926138e-06, 1.0926961e-07, -2.772859e-08, -4.7492586e-06, 1.7844712e-06, 8.040899e-08, -2.745329e-08, -3.8386715e-06, 1.854135e-06, 5.110077e-08, -2.6864837e-08, -2.8988977e-06, 1.9011702e-06, 2.16917e-08, -2.5975288e-08, -1.9413042e-06, 1.9254112e-06, -7.476121e-09, -2.4799975e-08, -9.772733e-07, 1.926959e-06, -3.6069117e-08, -2.335729e-08, -1.807226e-08, 1.9061755e-06, -6.3765945e-08, -2.1668402e-08, 9.252769e-07, 1.8636753e-06, -9.026101e-08, -1.9756987e-08, 1.8421199e-06, 1.800314e-06, -1.1526775e-07, -1.764889e-08, 2.7222877e-06, 1.717174e-06, -1.3852163e-07, -1.5371805e-08, 3.5562061e-06, 1.6155491e-06, -1.5978283e-07, -1.295492e-08, 4.3349964e-06, 1.4969248e-06, -1.788386e-07, -1.0428548e-08, 5.0505664e-06, 1.3629591e-06, -1.9550531e-07, -7.823766e-09, 5.695692e-06, 1.2154594e-06, -2.0963e-07, -5.172035e-09, 6.264085e-06, 1.0563596e-06, -2.2109177e-07, -2.504836e-09, 6.75045e-06, 8.8769553e-07, -2.2980251e-07, 1.4670004e-10, 7.150531e-06, 7.115797e-07, -2.3570743e-07, 2.7521438e-09, 7.4611416e-06, 5.301753e-07, -2.387852e-07, 5.282109e-09, 7.680183e-06, 3.456709e-07, -2.3904747e-07, 7.708576e-09, 7.806654e-06, 1.6025395e-07, -2.3653838e-07, 1.000519e-08, 7.840639e-06, -2.391398e-08, -2.3133336e-07, 1.2147542e-08, 7.783295e-06, -2.0472201e-07, -2.2353777e-07, 1.4113417e-08, 7.636812e-06, -3.8013349e-07, -2.1328523e-07, 1.5883016e-08, 7.40438e-06, -5.482083e-07, -2.0073556e-07, 1.7439138e-08, 7.090127e-06, -7.071237e-07, -1.8607247e-07, 1.876735e-08, 6.699061e-06, -8.5519366e-07, -1.6950105e-07, 1.985609e-08, 6.2369945e-06, -9.908856e-07, -1.5124509e-07, 2.0696767e-08, 5.7104644e-06, -1.1128363e-06, -1.315441e-07, 2.1283801e-08, 5.1266447e-06, -1.219864e-06, -1.1065032e-07, 2.1614644e-08, 4.4932526e-06, -1.3109797e-06, -8.882555e-08, 2.168976e-08, 3.8184494e-06, -1.385395e-06, -6.633802e-08, 2.1512554e-08, 3.1107395e-06, -1.4425282e-06, -4.3459114e-08, 2.1089306e-08, 2.3788657e-06, -1.4820073e-06, -2.046021e-08, 2.0429034e-08, 1.6317043e-06, -1.5036707e-06, 2.390464e-09, 1.9543348e-08, 8.781599e-07, -1.5075659e-06, 2.4830888e-08, 1.8446276e-08, 1.2706168e-07, -1.4939454e-06, 4.6608175e-08, 1.7154052e-08, -6.12937e-07, -1.4632601e-06, 6.748136e-08, 1.5684906e-08, -1.3334562e-06, -1.4161506e-06, 8.722395e-08, 1.4058801e-08, -2.0264818e-06, -1.3534374e-06, 1.0562636e-07, 1.229719e-08, -2.684452e-06, -1.2761074e-06, 1.2249802e-07, 1.0422732e-08, -3.3003373e-06, -1.1853006e-06, 1.3766926e-07, 8.459013e-09, -3.8677135e-06, -1.0822936e-06, 1.5099292e-07, 6.430259e-09, -4.3808245e-06, -9.68483e-07, 1.6234573e-07, 4.3610413e-09, -4.8346396e-06, -8.453671e-07, 1.7162925e-07, 2.2759892e-09, -5.2248984e-06, -7.145266e-07, 1.7877069e-07, 1.9950301e-10, -5.548147e-06, -5.776055e-07, 1.8372322e-07, -1.844525e-09, -5.801766e-06, -4.362903e-07, 1.8646618e-07, -3.832978e-09, -5.9839845e-06, -2.9229045e-07, 1.8700479e-07, -5.7437695e-09, -6.093889e-06, -1.4731768e-07, 1.8536974e-07, -7.556082e-09, -6.1314176e-06, -3.0663436e-09, 1.8161633e-07, -9.250585e-09, -6.097348e-06, 1.3880587e-07, 1.7582347e-07, -1.08096385e-08, -5.9932718e-06, 2.766966e-07, 1.6809237e-07, -1.2217463e-08, -5.8215664e-06, 4.090764e-07, 1.5854495e-07, -1.3460292e-08, -5.585351e-06, 5.3450515e-07, 1.4732214e-07, -1.4526505e-08, -5.28844e-06, 6.5164744e-07, 1.345819e-07, -1.5406716e-08, -4.935286e-06, 7.592859e-07, 1.2049708e-07, -1.6093848e-08, -4.5309184e-06, 8.563338e-07, 1.0525326e-07, -1.6583183e-08, -4.0808745e-06, 9.418451e-07, 8.904626e-08, -1.6872365e-08, -3.5911287e-06, 1.015023e-06, 7.2079835e-08, -1.69614e-08, -3.0680144e-06, 1.075227e-06, 5.4563067e-08, -1.6852606e-08, -2.518145e-06, 1.1219774e-06, 3.6707938e-08, -1.6550556e-08, -1.9483334e-06, 1.1549583e-06, 1.8726793e-08, -1.606198e-08, -1.3655091e-06, 1.1740184e-06, 8.2987467e-10, -1.5395658e-08, -7.766358e-07, 1.1791701e-06, -1.6777065e-08, -1.4562276e-08, -1.886312e-07, 1.1705865e-06, -3.3895077e-08, -1.3574279e-08, 3.9171306e-07, 1.1485972e-06, -5.0334197e-08, -1.2445691e-08, 9.578077e-07, 1.1136808e-06, -6.591551e-08, -1.1191929e-08, 1.5033388e-06, 1.066458e-06, -8.0473e-08, -9.829603e-09, 2.0223358e-06, 1.0076815e-06, -9.385532e-08, -8.376298e-09, 2.5092359e-06, 9.3822496e-07, -1.05927235e-07, -6.85036e-09, 2.95894e-06, 8.590712e-07, -1.1657094e-07, -5.270668e-09, 3.366866e-06, 7.712987e-07, -1.2568714e-07, -3.6564072e-09, 3.728991e-06, 6.760677e-07, -1.3319588e-07, -2.0268422e-09, 4.0418904e-06, 5.7460545e-07, -1.3903717e-07, -4.0109174e-10, 4.3027667e-06, 4.681907e-07, -1.4317129e-07, 1.2020895e-09, 4.5094707e-06, 3.581381e-07, -1.4557898e-07, 2.7645222e-09, 4.660517e-06, 2.457824e-07, -1.4626126e-07, 4.2688026e-09, 4.7550884e-06, 1.3246272e-07, -1.4523911e-07, 5.698492e-09, 4.7930366e-06, 1.9506862e-08, -1.4255292e-07, 7.0382895e-09, 4.7748695e-06, -9.178376e-08, -1.3826161e-07, 8.274192e-09, 4.7017375e-06, -2.0014883e-07, -1.3244174e-07, 9.393632e-09, 4.5754064e-06, -3.0438298e-07, -1.2518626e-07, 1.0385602e-08, 4.39823e-06, -4.0334885e-07, -1.1660318e-07, 1.1240753e-08, 4.17311e-06, -4.9598907e-07, -1.0681408e-07, 1.1951477e-08, 3.903455e-06, -5.8133725e-07, -9.595246e-08, 1.2511965e-08, 3.5931316e-06, -6.585275e-07, -8.4162e-08, 1.2918243e-08, 3.246413e-06, -7.268029e-07, -7.159472e-08, 1.3168191e-08, 2.8679215e-06, -7.8552245e-07, -5.8409096e-08, 1.3261532e-08, 2.4625701e-06, -8.3416637e-07, -4.4768104e-08, 1.3199808e-08, 2.0355008e-06, -8.723403e-07, -3.0837267e-08, 1.29863285e-08, 1.5920206e-06, -8.9977766e-07, -1.6782687e-08, 1.2626104e-08, 1.1375372e-06, -9.163406e-07, -2.7691178e-09, 1.2125762e-08, 6.7749596e-07, -9.220194e-07, 1.1041917e-08, 1.1493438e-08, 2.1731475e-07, -9.169306e-07, 2.4493941e-08, 1.0738662e-08, -2.3767731e-07, -9.0131334e-07, 3.7437257e-08, 9.872221e-09, -6.823005e-07, -8.755247e-07, 4.973056e-08, 8.906012e-09, -1.1115818e-06, -8.4003335e-07, 6.124243e-08, 7.852889e-09, -1.520809e-06, -7.954126e-07, 7.185271e-08, 6.7264976e-09, -1.9055809e-06, -7.423318e-07, 8.145366e-08, 5.5411027e-09, -2.2618533e-06, -6.8154696e-07, 8.995106e-08, 4.3114126e-09, -2.585979e-06, -6.1389073e-07, 9.726501e-08, 3.0524028e-09, -2.8747447e-06, -5.4026117e-07, 1.0333066e-07, 1.7791372e-09, -3.1253996e-06, -4.616106e-07, 1.0809872e-07, 5.065927e-10, -3.3356807e-06, -3.789335e-07, 1.115357e-07, -7.505129e-10, -3.5038295e-06, -2.9325426e-07, 1.13624104e-07, -1.9778867e-09, -3.628605e-06, -2.0561488e-07, 1.1436234e-07, -3.16182e-09, -3.709289e-06, -1.1706265e-07, 1.1376446e-07, -4.289335e-09, -3.745686e-06, -2.8637835e-08, 1.1185975e-07, -5.3483262e-09, -3.7381158e-06, 5.863815e-08, 1.08692134e-07, -6.3276815e-09, -3.687402e-06, 1.437743e-07, 1.0431943e-07, -7.2173987e-09, -3.5948542e-06, 2.2582097e-07, 9.8812414e-08, -8.00868e-09, -3.462244e-06, 3.0388017e-07, 9.225383e-08, -8.694013e-09, -3.2917767e-06, 3.771151e-07, 8.473719e-08, -9.267239e-09, -3.0860597e-06, 4.447588e-07, 7.6365545e-08, -9.723601e-09, -2.848064e-06, 5.061219e-07, 6.7250106e-08, -1.0059771e-08, -2.5810848e-06, 5.6059923e-07, 5.7508842e-08, -1.0273871e-08, -2.2886982e-06, 6.0767553e-07, 4.7264983e-08, -1.0365465e-08, -1.9747133e-06, 6.469297e-07, 3.664552e-08, -1.0335545e-08, -1.6431266e-06, 6.7803836e-07, 2.5779663e-08, -1.0186492e-08, -1.2980707e-06, 7.007778e-07, 1.479731e-08, -9.922023e-09, -9.4376543e-07, 7.1502484e-07, 3.827534e-09, -9.547135e-09, -5.8446665e-07, 7.2075676e-07, -7.002899e-09, -9.068013e-09, -2.2441691e-07, 7.180498e-07, -1.7570958e-08, -8.491949e-09, 1.3220347e-07, 7.0707654e-07, -2.7758706e-08, -7.827235e-09, 4.813239e-07, 6.8810243e-07, -3.7454587e-08, -7.0830475e-09, 8.190289e-07, 6.614809e-07, -4.65546e-08, -6.2693317e-09, 1.1416005e-06, 6.2764826e-07, -5.496339e-08, -5.3966707e-09, 1.445558e-06, 5.871168e-07, -6.25952e-08, -4.4761523e-09, 1.7276949e-06, 5.404678e-07, -6.937468e-08, -3.5192327e-09, 1.9851104e-06, 4.883437e-07, -7.5237644e-08, -2.537598e-09, 2.215239e-06, 4.3143942e-07, -8.013156e-08, -1.5430243e-09, 2.4158735e-06, 3.7049375e-07, -8.401601e-08, -5.472409e-10, 2.5851853e-06, 3.0627973e-07, -8.686292e-08, 4.3820567e-10, 2.7217388e-06, 2.395954e-07, -8.865671e-08, 1.4020818e-09, 2.824502e-06, 1.7125402e-07, -8.939425e-08, 2.3335915e-09, 2.8928507e-06, 1.02074345e-07, -8.908468e-08, 3.2224943e-09, 2.92657e-06, 3.2871213e-08, -8.774912e-08, 4.0592143e-09, 2.9258495e-06, -3.555395e-08, -8.54202e-08, 4.8349396e-09, 2.8912737e-06, -1.02422135e-07, -8.2141504e-08, 5.5417124e-09, 2.8238098e-06, -1.6698539e-07, -7.796689e-08, 6.172506e-09, 2.7247893e-06, -2.2853496e-07, -7.295968e-08, 6.7212906e-09, 2.5958864e-06, -2.8640886e-07, -6.719176e-08, 7.183087e-09, 2.4390934e-06, -3.3999873e-07, -6.074264e-08, 7.554006e-09, 2.2566924e-06, -3.8875592e-07, -5.3698376e-08, 7.831276e-09, 2.0512232e-06, -4.3219703e-07, -4.615046e-08, 8.013254e-09, 1.8254502e-06, -4.6990817e-07, -3.81947e-08, 8.0994305e-09, 1.582327e-06, -5.0154875e-07, -2.993001e-08, 8.09041e-09, 1.3249578e-06, -5.2685414e-07, -2.1457227e-08, 7.987892e-09, 1.0565604e-06, -5.456375e-07, -1.2877911e-08, 7.794628e-09, 7.804263e-07, -5.577906e-07, -4.2931516e-09, 7.514375e-09, 4.998811e-07, -5.6328366e-07, 4.1975903e-09, 7.151831e-09, 2.1824597e-07, -5.6216476e-07, 1.2497605e-08, 6.7125727e-09, -6.1200744e-08, -5.545574e-07, 2.0514012e-08, 6.2029675e-09, -3.352611e-07, -5.406583e-07, 2.8158766e-08, 5.630092e-09, -6.008529e-07, -5.207337e-07, 3.53496e-08, 5.0016364e-09, -8.5504377e-07, -4.9511505e-07, 4.201088e-08, 4.3258064e-09, -1.0950822e-06, -4.641942e-07, 4.807436e-08, 3.6112175e-09, -1.3184266e-06, -4.2841788e-07, 5.3479866e-08, 2.86679e-09, -1.5227712e-06, -3.8828145e-07, 5.817584e-08, 2.1016404e-09, -1.7060687e-06, -3.4432253e-07, 6.21198e-08, 1.3249726e-09, -1.8665498e-06, -2.971139e-07, 6.527869e-08, 5.459693e-10, -2.002739e-06, -2.4725642e-07, 6.762909e-08, -2.2631316e-10, -2.1134663e-06, -1.9537156e-07, 6.915731e-08, -9.83048e-10, -2.1978763e-06, -1.4209381e-07, 6.9859446e-08, -1.715736e-09, -2.2554327e-06, -8.806321e-08, 6.974118e-08, -2.4162987e-09, -2.2859185e-06, -3.391776e-08, 6.8817634e-08, -3.0771647e-09, -2.2894344e-06, 1.9713866e-08, 6.711297e-08, -3.6913492e-09, -2.266391e-06, 7.221948e-08, 6.465999e-08, -4.2525237e-09, -2.2174995e-06, 1.2301017e-07, 6.149963e-08, -4.7550803e-09, -2.1437586e-06, 1.7152672e-07, 5.76803e-08, -5.1941833e-09, -2.046438e-06, 2.1724563e-07, 5.3257242e-08, -5.565812e-09, -1.927059e-06, 2.5968453e-07, 4.8291767e-08, -5.8667937e-09, -1.7873724e-06, 2.9840706e-07, 4.2850427e-08, -6.0948278e-09, -1.6293353e-06, 3.3302726e-07, 3.7004174e-08, -6.248496e-09, -1.4550841e-06, 3.6321305e-07, 3.0827458e-08, -6.327264e-09, -1.2669072e-06, 3.8868924e-07, 2.4397309e-08, -6.331474e-09, -1.0672161e-06, 4.092398e-07, 1.7792399e-08, -6.2623253e-09, -8.585148e-07, 4.247093e-07, 1.1092104e-08, -6.121847e-09, -6.4336996e-07, 4.3500376e-07, 4.3755817e-09, -5.912858e-09, -4.2437983e-07, 4.4009064e-07, -2.2791529e-09, -5.6389258e-09, -2.0414359e-07, 4.3999825e-07, -8.796104e-09, -5.304307e-09, 1.47686166e-08, 4.3481432e-07, -1.5102144e-08, -4.913892e-09, 2.2984501e-07, 4.2468412e-07, -2.1127807e-08, -4.473133e-09, 4.3866027e-07, 4.098077e-07, -2.6808044e-08, -3.9879753e-09, 6.389021e-07, 3.9043675e-07, -3.208288e-08, -3.4647774e-09, 8.2839625e-07, 3.6687072e-07, -3.6898054e-08, -2.9102325e-09, 1.0051291e-06, 3.3945258e-07, -4.1205517e-08, -2.3312843e-09, 1.1672687e-06, 3.0856424e-07, -4.496391e-08, -1.7350429e-09, 1.3131826e-06, 2.7462127e-07, -4.8138922e-08, -1.128699e-09, 1.4414532e-06, 2.3806776e-07, -5.070357e-08, -5.194406e-10, 1.5508913e-06, 1.993705e-07, -5.2638377e-08, 8.563136e-11, 1.6405454e-06, 1.5901331e-07, -5.39315e-08, 6.795831e-10, 1.7097088e-06, 1.1749112e-07, -5.457871e-08, 1.2557257e-09, 1.7579241e-06, 7.530406e-08, -5.4583328e-08, 1.8076884e-09, 1.7849839e-06, 3.2951583e-08, -5.3956057e-08, 2.3294868e-09, 1.790929e-06, -9.073299e-09, -5.2714736e-08, 2.815586e-09, 1.7760442e-06, -5.028963e-08, -5.0884015e-08, 3.260957e-09, 1.7408503e-06, -9.023385e-08, -4.849495e-08, 3.6611263e-09, 1.686095e-06, -1.284649e-07, -4.5584542e-08, 4.0122186e-09, 1.6127392e-06, -1.6456893e-07, -4.2195207e-08, 4.3109916e-09, 1.5219435e-06, -1.9816363e-07, -3.8374196e-08, 4.5548623e-09};
	localparam real hb[0:3999] = {0.024986578, 0.000116877105, -3.896343e-05, -2.2712003e-07, 0.024869869, 0.0003495672, -3.6725352e-05, -6.683011e-07, 0.02463752, 0.00057908345, -3.2282736e-05, -1.071189e-06, 0.02429164, 0.00080335606, -2.5699466e-05, -1.4122909e-06, 0.023835355, 0.0010203768, -1.7068134e-05, -1.6701244e-06, 0.023272775, 0.0012282217, -6.508329e-06, -1.825436e-06, 0.02260895, 0.0014250721, 5.835373e-06, -1.8613864e-06, 0.021849804, 0.0016092348, 1.979567e-05, -1.7637041e-06, 0.021002075, 0.0017791594, 3.5185032e-05, -1.5208042e-06, 0.020073237, 0.0019334549, 5.1798383e-05, -1.1238726e-06, 0.019071415, 0.0020709035, 6.941594e-05, -5.669145e-07, 0.018005302, 0.0021904726, 8.7806206e-05, 1.5323168e-07, 0.016884053, 0.0022913238, 0.000106729, 1.0369153e-06, 0.015717195, 0.0023728213, 0.00012593858, 2.0817276e-06, 0.014514523, 0.0024345345, 0.00014518676, 3.2825897e-06, 0.01328599, 0.0024762424, 0.000164226, 4.6318687e-06, 0.012041612, 0.0024979326, 0.00018281244, 6.119525e-06, 0.010791358, 0.0024997983, 0.00020070883, 7.733287e-06, 0.009545049, 0.0024822343, 0.00021768737, 9.458844e-06, 0.008312262, 0.0024458296, 0.00023353235, 1.1280068e-05, 0.0071022296, 0.0023913574, 0.00024804258, 1.31792485e-05, 0.0059237573, 0.0023197657, 0.0002610337, 1.5137347e-05, 0.004785133, 0.0022321627, 0.00027234023, 1.7134254e-05, 0.003694055, 0.002129803, 0.00028181716, 1.9149073e-05, 0.0026575602, 0.0020140712, 0.0002893417, 2.116038e-05, 0.0016819648, 0.0018864649, 0.00029481426, 2.3146522e-05, 0.0007728115, 0.0017485761, 0.00029815955, 2.5085883e-05, -6.517271e-05, 0.0016020724, 0.00029932705, 2.6957157e-05, -0.0008281093, 0.0014486772, 0.0002982914, 2.8739623e-05, -0.0015129913, 0.0012901495, 0.00029505236, 3.0413386e-05, -0.002117696, 0.0011282647, 0.0002896347, 3.195963e-05, -0.0026409882, 0.00096479343, 0.0002820874, 3.3360822e-05, -0.003082513, 0.00080148317, 0.00027248287, 3.4600955e-05, -0.0034427792, 0.00064003846, 0.000260916, 3.5665686e-05, -0.0037231334, 0.0004821034, 0.00024750258, 3.6542533e-05, -0.003925726, 0.00032924407, 0.00023237792, 3.7221005e-05, -0.004053466, 0.00018293266, 0.00021569492, 3.76927e-05, -0.0041099745, 4.453296e-05, 0.00019762217, 3.79514e-05, -0.0040995227, -8.471297e-05, 0.00017834186, 3.7993144e-05, -0.0040269704, -0.00020369625, 0.00015804752, 3.7816237e-05, -0.0038976963, -0.00031145103, 0.00013694167, 3.742127e-05, -0.0037175252, -0.00040716256, 0.00011523339, 3.6811085e-05, -0.0034926496, -0.0004901733, 9.3135954e-05, 3.599074e-05, -0.0032295508, -0.00055998715, 7.086427e-05, 3.4967423e-05, -0.002934917, -0.0006162719, 4.8632493e-05, 3.3750366e-05, -0.0026155617, -0.0006588598, 2.6651622e-05, 3.235072e-05, -0.0022783414, -0.0006877456, 5.1271536e-06, 3.0781408e-05, -0.0019300748, -0.00070308376, -1.5743133e-05, 2.9056979e-05, -0.0015774649, -0.0007051833, -3.577129e-05, 2.7193415e-05, -0.0012270228, -0.00069450086, -5.4781158e-05, 2.5207955e-05, -0.00088499615, -0.00067163265, -7.261017e-05, 2.311889e-05, -0.00055730145, -0.0006373044, -8.911096e-05, 2.0945343e-05, -0.0002494623, -0.00059236056, -0.00010415277, 1.8707058e-05, 3.3447053e-05, -0.00053775206, -0.00011762269, 1.6424181e-05, 0.00028685166, -0.00047452268, -0.00012942658, 1.4117025e-05, 0.0005067189, -0.00040379557, -0.0001394899, 1.1805854e-05, 0.00068959437, -0.00032675808, -0.00014775814, 9.510665e-06, 0.0008326304, -0.00024464677, -0.00015419716, 7.2509692e-06, 0.0009336064, -0.00015873181, -0.00015879319, 5.0455933e-06, 0.0009909424, -7.03015e-05, -0.0001615527, 2.9124817e-06, 0.0010037036, 1.9353303e-05, -0.00016250192, 8.6851696e-07, 0.000971598, 0.00010895448, -0.00016168621, -1.0706473e-06, 0.00089496677, 0.00019725144, -0.00015916926, -2.890736e-06, 0.0007747661, 0.0002830354, -0.00015503199, -4.578985e-06, 0.0006125435, 0.0003651528, -0.0001493714, -6.1242554e-06, 0.00041040673, 0.00044251818, -0.00014229909, -7.517124e-06, 0.00017098685, 0.0005141254, -0.00013393987, -8.749958e-06, -0.000102604055, 0.0005790583, -0.00012442996, -9.816967e-06, -0.00040682033, 0.00063650013, -0.00011391535, -1.0714228e-05, -0.0007377343, 0.00068574096, -0.000102549915, -1.1439698e-05, -0.0010910918, 0.00072618475, -9.049353e-05, -1.1993197e-05, -0.0014623696, 0.0007573539, -7.791015e-05, -1.237638e-05, -0.0018468365, 0.0007788933, -6.496585e-05, -1.2592673e-05, -0.002239615, 0.0007905721, -5.1826923e-05, -1.2647208e-05, -0.0026357428, 0.0007922844, -3.8657945e-05, -1.2546729e-05, -0.0030302363, 0.00078404846, -2.5619947e-05, -1.22994825e-05, -0.0034181513, 0.0007660045, -1.2868641e-05, -1.1915097e-05, -0.0037946438, 0.0007384107, -5.527264e-07, -1.1404446e-05, -0.0041550267, 0.00070163846, 1.1187671e-05, -1.0779499e-05, -0.0044948263, 0.000656166, 2.2222448e-05, -1.0053163e-05, -0.004809833, 0.00060257106, 3.2432832e-05, -9.239121e-06, -0.005096149, 0.0005415224, 4.1712527e-05, -8.351654e-06, -0.0053502326, 0.00047377063, 4.9968694e-05, -7.4054738e-06, -0.0055689337, 0.0004001377, 5.7122783e-05, -6.415538e-06, -0.005749531, 0.00032150644, 6.311115e-05, -5.3968797e-06, -0.005889757, 0.00023880896, 6.788551e-05, -4.3644327e-06, -0.005987819, 0.00015301503, 7.1413204e-05, -3.33286e-06, -0.0060424167, 6.5120075e-05, 7.367729e-05, -2.3163923e-06, -0.0060527516, -2.3866987e-05, 7.467643e-05, -1.3286729e-06, -0.006018531, -0.00011293571, 7.442458e-05, -3.8261123e-07, -0.0059399647, -0.00020108608, 7.295059e-05, 5.097503e-07, -0.005817757, -0.00028734, 7.029756e-05, 1.3373586e-06, -0.0056530945, -0.00037075247, 6.652203e-05, 2.0902578e-06, -0.005447625, -0.00045042214, 6.169313e-05, 2.759682e-06, -0.0052034347, -0.00052550115, 5.589148e-05, 3.3381343e-06, -0.004923017, -0.00059520424, 4.9208058e-05, 3.819447e-06, -0.004609243, -0.00065881707, 4.1742933e-05, 4.198827e-06, -0.0042653196, -0.0007157032, 3.3603916e-05, 4.472884e-06, -0.003894752, -0.0007653107, 2.4905143e-05, 4.639643e-06, -0.0035012984, -0.0008071772, 1.5765636e-05, 4.698537e-06, -0.003088926, -0.0008409337, 6.307793e-06, 4.6503856e-06, -0.0026617618, -0.0008663077, -3.3441117e-06, 4.4973604e-06, -0.0022240446, -0.00088312494, -1.3065424e-05, 4.2429283e-06, -0.0017800763, -0.0008913099, -2.2732595e-05, 3.8917874e-06, -0.0013341709, -0.000890885, -3.2224616e-05, 3.4497868e-06, -0.0008906079, -0.00088196935, -4.142441e-05, 2.9238345e-06, -0.0004535831, -0.00086477544, -5.0220144e-05, 2.321794e-06, -2.7163756e-05, -0.00083960575, -5.850646e-05, 1.652374e-06, 0.00038475564, -0.0008068475, -6.618562e-05, 9.250065e-07, 0.0007784943, -0.0007669673, -7.316853e-05, 1.497222e-07, 0.0011506232, -0.00072050426, -7.937563e-05, -6.629815e-07, 0.0014979994, -0.000668063, -8.473774e-05, -1.5022744e-06, 0.0018177973, -0.0006103056, -8.919661e-05, -2.3571292e-06, 0.0021075346, -0.000547943, -9.270552e-05, -3.2164576e-06, 0.002365095, -0.00048172637, -9.522962e-05, -4.069244e-06, 0.002588746, -0.00041243774, -9.674611e-05, -4.9046766e-06, 0.0027771518, -0.00034088065, -9.7244396e-05, -5.7122747e-06, 0.0029293816, -0.00026787055, -9.672597e-05, -6.482007e-06, 0.0030449138, -0.00019422543, -9.520421e-05, -7.204406e-06, 0.0031236338, -0.00012075634, -9.270407e-05, -7.870673e-06, 0.0031658295, -4.8258335e-05, -8.926157e-05, -8.472772e-06, 0.0031721801, 2.2498389e-05, -8.492326e-05, -9.003513e-06, 0.003143742, 9.077683e-05, -7.974546e-05, -9.4566285e-06, 0.0030819303, 0.00015588106, -7.379349e-05, -9.826832e-06, 0.0029884963, 0.00021716346, -6.714076e-05, -1.0109866e-05, 0.0028655012, 0.00027403128, -5.9867805e-05, -1.030254e-05, 0.0027152882, 0.00032595254, -5.206122e-05, -1.0402753e-05, 0.0025404498, 0.000372461, -4.3812594e-05, -1.04095e-05, 0.0023437948, 0.0004131604, -3.5217337e-05, -1.032287e-05, 0.0021283112, 0.0004477277, -2.6373558e-05, -1.0144035e-05, 0.0018971302, 0.0004759157, -1.738085e-05, -9.875211e-06, 0.0016534871, 0.0004975543, -8.339134e-06, -9.5196265e-06, 0.001400683, 0.0005125514, 6.5249236e-07, -9.081469e-06, 0.0011420455, 0.00052089227, 9.4969e-06, -8.565822e-06, 0.00088089047, 0.00052263855, 1.810001e-05, -7.978593e-06, 0.00062048424, 0.0005179262, 2.6371838e-05, -7.3264337e-06, 0.00036400717, 0.0005069625, 3.422745e-05, -6.6166567e-06, 0.00011451893, 0.00049002253, 4.1587886e-05, -5.8571363e-06, -0.0001250745, 0.0004674449, 4.8380953e-05, -5.0562144e-06, -0.0003520511, 0.00043962628, 5.4541957e-05, -4.222595e-06, -0.0005639008, 0.00040701643, 6.0014332e-05, -3.365242e-06, -0.00075835024, 0.0003701115, 6.475016e-05, -2.4932692e-06, -0.0009333844, 0.00032944788, 6.871057e-05, -1.6158366e-06, -0.0010872651, 0.00028559507, 7.186606e-05, -7.4204394e-07, -0.0012185457, 0.00023914858, 7.419667e-05, 1.1917229e-07, -0.0013260824, 0.00019072261, 7.5692085e-05, 9.591386e-07, -0.0014090413, 0.00014094257, 7.635154e-05, 1.7695393e-06, -0.0014669029, 9.043767e-05, 7.6183744e-05, 2.5425059e-06, -0.0014994614, 3.9833558e-05, 7.5206575e-05, 3.2706998e-06, -0.0015068215, -1.0254878e-05, 7.344675e-05, 3.9473884e-06, -0.0014893912, -5.9230428e-05, 7.093935e-05, 4.566511e-06, -0.0014478713, -0.00010652019, 6.772732e-05, 5.122739e-06, -0.0013832418, -0.00015158176, 6.386082e-05, 5.6115227e-06, -0.0012967449, -0.00019390904, 5.93965e-05, 6.0291327e-06, -0.0011898658, -0.00023303744, 5.4396824e-05, 6.372689e-06, -0.0010643104, -0.00026854855, 4.8929178e-05, 6.6401776e-06, -0.0009219817, -0.0003000742, 4.3065043e-05, 6.830463e-06, -0.0007649533, -0.00032729987, 3.6879126e-05, 6.943284e-06, -0.00059544214, -0.00034996742, 3.0448418e-05, 6.9792427e-06, -0.00041577968, -0.00036787707, 2.3851286e-05, 6.9397847e-06, -0.0002283824, -0.00038088873, 1.716655e-05, 6.827166e-06, -3.5721743e-05, -0.0003889226, 1.0472569e-05, 6.6444177e-06, 0.00015970602, -0.00039195913, 3.84635e-06, 6.3952925e-06, 0.0003554097, -0.00039003804, -2.637314e-06, 6.0842167e-06, 0.0005489325, -0.000383257, -8.906665e-06, 5.7162215e-06, 0.0007378806, -0.00037176942, -1.4893752e-05, 5.2968808e-06, 0.00091995014, -0.0003557817, -2.0535148e-05, 4.8322336e-06, 0.0010929531, -0.00033554994, -2.5772597e-05, 4.328711e-06, 0.0012548412, -0.00031137612, -3.0553598e-05, 3.7930529e-06, 0.0014037276, -0.00028360382, -3.483191e-05, 3.2322278e-06, 0.0015379067, -0.00025261342, -3.8567974e-05, 2.653347e-06, 0.0016558714, -0.00021881713, -4.172925e-05, 2.0635835e-06, 0.0017563275, -0.00018265363, -4.4290467e-05, 1.4700853e-06, 0.0018382053, -0.0001445825, -4.6233796e-05, 8.798973e-07, 0.0019006693, -0.00010507852, -4.7548918e-05, 2.9988044e-07, 0.001943124, -6.462584e-05, -4.8233018e-05, -2.63363e-07, 0.0019652168, -2.3712253e-05, -4.829067e-05, -8.035608e-07, 0.001966839, 1.7176591e-05, -4.7733673e-05, -1.3148367e-06, 0.0019481225, 5.7562815e-05, -4.6580783e-05, -1.7917708e-06, 0.001909436, 9.6981734e-05, -4.4857356e-05, -2.229454e-06, 0.0018513753, 0.00013498706, -4.2594966e-05, -2.6235343e-06, 0.0017747541, 0.00017115581, -3.983091e-05, -2.9702587e-06, 0.0016805907, 0.00020509283, -3.6607682e-05, -3.2665032e-06, 0.0015700932, 0.00023643493, -3.2972388e-05, -3.5097996e-06, 0.0014446424, 0.00026485464, -2.8976121e-05, -3.6983504e-06, 0.0013057735, 0.00029006338, -2.4673294e-05, -3.8310386e-06, 0.0011551554, 0.0003118142, -2.012095e-05, -3.907428e-06, 0.0009945696, 0.00032990403, -1.537806e-05, -3.9277547e-06, 0.00082588807, 0.00034417518, -1.0504799e-05, -3.892914e-06, 0.0006510498, 0.0003545167, -5.5618216e-06, -3.8044357e-06, 0.00047203756, 0.0003608646, -6.095561e-07, -3.6644583e-06, 0.0002908543, 0.0003632021, 4.2925003e-06, -3.4756895e-06, 0.00010949978, 0.0003615589, 9.086454e-06, -3.2413664e-06, -7.005265e-05, 0.00035601013, 1.3716667e-05, -2.9652074e-06, -0.00024587815, 0.00034667485, 1.8130359e-05, -2.6513612e-06, -0.000416122, 0.00033371375, 2.2278178e-05, -2.3043497e-06, -0.00057901966, 0.00031732683, 2.6114716e-05, -1.929009e-06, -0.0007329159, 0.00029775038, 2.959897e-05, -1.5304275e-06, -0.00087628193, 0.00027525355, 3.269475e-05, -1.1138819e-06, -0.0010077311, 0.00025013494, 3.5371e-05, -6.847718e-07, -0.0011260324, 0.00022271842, 3.760211e-05, -2.4855487e-07, -0.0012301225, 0.00019334916, 3.936808e-05, 1.893183e-07, -0.001319115, 0.00016238925, 4.0654697e-05, 6.234677e-07, -0.0013923077, 0.0001302132, 4.1453575e-05, 1.0486458e-06, -0.0014491879, 9.720347e-05, 4.1762174e-05, 1.4597965e-06, -0.0014894352, 6.374589e-05, 4.1583724e-05, 1.8521115e-06, -0.0015129221, 3.0225176e-05, 4.092709e-05, 2.221082e-06, -0.0015197119, -2.9794865e-06, 3.980659e-05, 2.5625463e-06, -0.0015100557, -3.5498742e-05, 3.8241713e-05, 2.8727338e-06, -0.0014843857, -6.697716e-05, 3.6256835e-05, 3.1483007e-06, -0.0014433075, -9.707708e-05, 3.388084e-05, 3.386364e-06, -0.0013875904, -0.00012548224, 3.1146705e-05, 3.584526e-06, -0.0013181557, -0.00015190107, 2.8091063e-05, 3.740896e-06, -0.0012360639, -0.00017606962, 2.4753714e-05, 3.854103e-06, -0.0011424997, -0.00019775413, 2.1177106e-05, 3.9233023e-06, -0.0010387572, -0.00021675328, 1.74058e-05, 3.9481793e-06, -0.0009262218, -0.00023289995, 1.3485926e-05, 3.928943e-06, -0.0008063545, -0.00024606255, 9.464609e-06, 3.866315e-06, -0.0006806726, -0.00025614596, 5.3894196e-06, 3.7615139e-06, -0.0005507317, -0.00026309196, 1.3078055e-06, 3.6162312e-06, -0.00041810746, -0.00026687945, -2.7334515e-06, 3.4326067e-06, -0.00028437664, -0.00026752386, -6.688769e-06, 3.2131943e-06, -0.00015109948, -0.0002650765, -1.0514272e-05, 2.9609264e-06, -1.9801768e-05, -0.00025962334, -1.4168271e-05, 2.6790735e-06, 0.00010804198, -0.00025128332, -1.7611716e-05, 2.3712018e-06, 0.00023102465, -0.00024020665, -2.0808595e-05, 2.041126e-06, 0.0003478215, -0.00022657229, -2.3726312e-05, 1.6928611e-06, 0.000457204, -0.0002105856, -2.6336e-05, 1.3305736e-06, 0.00055805227, -0.0001924754, -2.86128e-05, 9.585298e-07, 0.0006493661, -0.00017249103, -3.053608e-05, 5.8104513e-07, 0.0007302744, -0.00015089898, -3.2089603e-05, 2.0243363e-07, 0.00080004294, -0.0001279797, -3.3261647e-05, -1.7304232e-07, 0.00085808046, -0.00010402399, -3.4045068e-05, -5.412203e-07, 0.000903943, -7.932951e-05, -3.4437293e-05, -8.9808447e-07, 0.0009373362, -5.4197226e-05, -3.4440294e-05, -1.2398096e-06, 0.00095811655, -2.8927887e-05, -3.4060486e-05, -1.5628023e-06, 0.00096629, -3.8185226e-06, -3.3308566e-05, -1.8637385e-06, 0.0009620094, 2.0840904e-05, -3.219934e-05, -2.139598e-06, 0.0009455702, 4.477073e-05, -3.075146e-05, -2.3876942e-06, 0.0009174042, 6.770467e-05, -2.8987177e-05, -2.6056998e-06, 0.00087807275, 8.939263e-05, -2.6931988e-05, -2.7916674e-06, 0.00082825747, 0.00010960339, -2.461432e-05, -2.9440466e-06, 0.0007687504, 0.00012812686, -2.2065136e-05, -3.0616948e-06, 0.0007004428, 0.00014477625, -1.9317536e-05, -3.1438838e-06, 0.0006243134, 0.00015938978, -1.6406348e-05, -3.1903023e-06, 0.000541415, 0.00017183211, -1.33676895e-05, -3.2010514e-06, 0.0004528613, 0.00018199554, -1.0238536e-05, -3.1766376e-06, 0.00035981278, 0.00018980069, -7.0562724e-06, -3.1179597e-06, 0.00026346243, 0.00019519699, -3.8582616e-06, -3.0262931e-06, 0.00016502131, 0.00019816274, -6.8140974e-07, -2.9032674e-06, 6.570411e-05, 0.00019870495, 2.4382505e-06, -2.7508431e-06, -3.3284992e-05, 0.00019685866, 5.465961e-06, -2.5712827e-06, -0.0001307662, 0.00019268612, 8.368619e-06, -2.3671205e-06, -0.00022559743, 0.0001862756, 1.111513e-05, -2.1411277e-06, -0.0003166869, 0.00017773996, 1.3676734e-05, -1.896278e-06, -0.00040300505, 0.00016721482, 1.6027298e-05, -1.635709e-06, -0.00048359542, 0.00015485672, 1.814357e-05, -1.3626835e-06, -0.0005575847, 0.00014084089, 2.0005407e-05, -1.0805502e-06, -0.00062419113, 0.00012535887, 2.1595948e-05, -7.927032e-07, -0.0006827326, 0.000108616085, 2.2901751e-05, -5.025426e-07, -0.0007326324, 9.082921e-05, 2.3912902e-05, -2.1343516e-07, -0.0007734245, 7.222342e-05, 2.4623056e-05, 7.132415e-08, -0.00080475706, 5.3029675e-05, 2.502946e-05, 3.4854867e-07, -0.0008263945, 3.3481938e-05, 2.513292e-05, 6.1519495e-07, -0.0008382184, 1.3814398e-05, 2.4937726e-05, 8.6839543e-07, -0.00084022695, -5.7412394e-06, 2.445156e-05, 1.1054885e-06, -0.000832533, -2.4958403e-05, 2.3685325e-05, 1.3240457e-06, -0.0008153609, -4.36182e-05, 2.2652985e-05, 1.5218957e-06, -0.00078904204, -6.151183e-05, 2.1371345e-05, 1.6971446e-06, -0.0007540092, -7.844284e-05, 1.98598e-05, 1.8481938e-06, -0.0007107897, -9.4229166e-05, 1.8140086e-05, 1.973753e-06, -0.0006599982, -0.00010870506, 1.6235963e-05, 2.072849e-06, -0.0006023276, -0.00012172271, 1.4172929e-05, 2.1448332e-06, -0.0005385399, -0.00013315363, 1.197788e-05, 2.189382e-06, -0.0004694564, -0.0001428899, 9.678783e-06, 2.2064958e-06, -0.00039594696, -0.000150845, 7.3043298e-06, 2.1964927e-06, -0.0003189192, -0.00015695447, 4.8835964e-06, 2.16e-06, -0.00023930735, -0.00016117636, 2.4456945e-06, 2.0979417e-06, -0.000158061, -0.00016349126, 1.9438557e-08, 2.0115217e-06, -7.613381e-05, -0.00016390221, -2.3669863e-06, 1.9022065e-06, 5.5276073e-06, -0.00016243423, -4.6863383e-06, 1.7717024e-06, 8.599451e-05, -0.00015913373, -6.91262e-06, 1.6219325e-06, 0.00016436652, -0.00015406757, -9.021357e-06, 1.4550101e-06, 0.0002397816, -0.000147322, -1.09898565e-05, 1.2732113e-06, 0.00031142536, -0.00013900126, -1.2797443e-05, 1.0789458e-06, 0.00037853981, -0.00012922616, -1.4425657e-05, 8.7472654e-07, 0.0004404311, -0.000118132346, -1.585844e-05, 6.631388e-07, 0.0004964765, -0.000105868516, -1.7082273e-05, 4.4680903e-07, 0.0005461306, -9.259446e-05, -1.8086295e-05, 2.2837375e-07, 0.0005889301, -7.847905e-05, -1.8862385e-05, 1.0448686e-08, 0.00062449806, -6.369811e-05, -1.94052e-05, -2.0440125e-07, 0.00065254676, -4.84323e-05, -1.9712208e-05, -4.1369077e-07, 0.0006728795, -3.2864893e-05, -1.9783653e-05, -6.150418e-07, 0.0006853914, -1.7179666e-05, -1.9622514e-05, -8.062092e-07, 0.00069006934, -1.5587267e-06, -1.9234425e-05, -9.851045e-07, 0.00068699016, 1.3819545e-05, -1.8627563e-05, -1.1498179e-06, 0.0006763186, 2.8782508e-05, -1.7812508e-05, -1.2986367e-06, 0.00065830396, 4.316516e-05, -1.6802087e-05, -1.4300626e-06, 0.0006332757, 5.6811925e-05, -1.5611182e-05, -1.5428252e-06, 0.0006016385, 6.957828e-05, -1.4256523e-05, -1.6358925e-06, 0.000563866, 8.1332255e-05, -1.2756469e-05, -1.7084797e-06, 0.00052049453, 9.195575e-05, -1.1130761e-05, -1.7600535e-06, 0.00047211576, 0.00010134568, -9.4002735e-06, -1.7903343e-06, 0.00041936894, 0.00010941489, -7.5867533e-06, -1.7992952e-06, 0.00036293277, 0.000116092924, -5.712553e-06, -1.7871583e-06, 0.00030351683, 0.00012132655, -3.8003616e-06, -1.7543875e-06, 0.00024185305, 0.00012508009, -1.8729359e-06, -1.7016795e-06, 0.00017868665, 0.00012733552, 4.716473e-08, -1.6299514e-06, 0.00011476754, 0.00012809242, 1.9378356e-06, -1.540327e-06, 5.0841467e-05, 0.0001273677, 3.7776758e-06, -1.43412e-06, -1.2358492e-05, 0.00012519505, 5.5462247e-06, -1.3128151e-06, -7.412017e-05, 0.000121624274, 7.224183e-06, -1.1780489e-06, -0.0001337602, 0.00011672055, 8.793616e-06, -1.0315878e-06, -0.00019063136, 0.00011056328, 1.0238141e-05, -8.753053e-07, -0.00024412952, 0.00010324503, 1.154309e-05, -7.1115886e-07, -0.00029369982, 9.487021e-05, 1.269565e-05, -5.4116543e-07, -0.00033884228, 8.555365e-05, 1.3684982e-05, -3.673775e-07, -0.00037911665, 7.541913e-05, 1.4502314e-05, -1.918583e-07, -0.00041414646, 6.459776e-05, 1.5141006e-05, -1.6657985e-08, -0.00044362227, 5.322641e-05, 1.5596595e-05, 1.5621004e-07, -0.00046730423, 4.1445935e-05, 1.5866808e-05, 3.2479178e-07, -0.00048502345, 2.9399558e-05, 1.5951551e-05, 4.872143e-07, -0.000496683, 1.7231143e-05, 1.5852878e-05, 6.417063e-07, -0.00050225767, 5.0835165e-06, 1.5574926e-05, 7.866165e-07, -0.000501793, -6.9031535e-06, 1.5123837e-05, 9.204313e-07, -0.00049540366, -1.8592944e-05, 1.4507653e-05, 1.0417896e-06, -0.00048327097, -2.985567e-05, 1.37361885e-05, 1.1494964e-06, -0.00046563946, -4.0568302e-05, 1.2820891e-05, 1.2425335e-06, -0.00044281324, -5.061626e-05, 1.17746795e-05, 1.3200689e-06, -0.00041515133, -5.989461e-05, 1.0611769e-05, 1.3814628e-06, -0.00038306252, -6.830909e-05, 9.347489e-06, 1.4262722e-06, -0.00034699994, -7.5777054e-05, 7.998085e-06, 1.4542526e-06, -0.00030745493, -8.22282e-05, 6.580511e-06, 1.4653576e-06, -0.0002649508, -8.760522e-05, 5.1122324e-06, 1.4597363e-06, -0.00022003613, -9.186418e-05, 3.6110046e-06, 1.437728e-06, -0.00017327811, -9.4974865e-05, 2.0946684e-06, 1.3998554e-06, -0.00012525555, -9.692086e-05, 5.8094145e-07, 1.3468156e-06, -7.655202e-05, -9.769953e-05, -9.127852e-07, 1.2794687e-06, -2.7749007e-05, -9.732179e-05, -2.3696427e-06, 1.198826e-06, 2.058078e-05, -9.581178e-05, -3.7734703e-06, 1.1060347e-06, 6.7879904e-05, -9.320637e-05, -5.1089905e-06, 1.0023633e-06, 0.000113612405, -8.955446e-05, -6.3619723e-06, 8.8918443e-07, 0.00015726963, -8.491628e-05, -7.5193757e-06, 7.6795754e-07, 0.00019837571, -7.9362464e-05, -8.569485e-06, 6.402103e-07, 0.00023649246, -7.2973075e-05, -9.502019e-06, 5.075201e-07, 0.00027122386, -6.5836495e-05, -1.0308231e-05, 3.7149482e-07, 0.00030221997, -5.8048292e-05, -1.0980981e-05, 2.3375374e-07, 0.0003291801, -4.970997e-05, -1.1514789e-05, 9.590874e-08, 0.0003518556, -4.09277e-05, -1.1905875e-05, -4.045425e-08, 0.0003700517, -3.1811025e-05, -1.2152172e-05, -1.7379317e-07, 0.0003836291, -2.247151e-05, -1.2253321e-05, -3.026269e-07, 0.00039250444, -1.3021434e-05, -1.2210649e-05, -4.2555126e-07, 0.00039665043, -3.5724718e-06, -1.2027122e-05, -5.4125417e-07, 0.00039609513, 5.7655866e-06, -1.1707282e-05, -6.48529e-07, 0.00039092085, 1.488608e-05, -1.1257177e-05, -7.46287e-07, 0.00038126216, 2.3686656e-05, -1.06842535e-05, -8.3356764e-07, 0.00036730347, 3.2070388e-05, -9.997255e-06, -9.095478e-07, 0.00034927618, 3.99468e-05, -9.206096e-06, -9.735488e-07, 0.00032745497, 4.7232814e-05, -8.32173e-06, -1.0250419e-06, 0.00030215413, 5.3853582e-05, -7.3560022e-06, -1.0636519e-06, 0.00027372318, 5.9743223e-05, -6.3214984e-06, -1.0891589e-06, 0.00024254216, 6.484542e-05, -5.231389e-06, -1.1014981e-06, 0.00020901674, 6.911395e-05, -4.0992645e-06, -1.1007583e-06, 0.00017357318, 7.2512994e-05, -2.9389716e-06, -1.0871773e-06, 0.00013665296, 7.501741e-05, -1.7644494e-06, -1.0611384e-06, 9.87074e-05, 7.6612865e-05, -5.895656e-07, -1.0231615e-06, 6.0192346e-05, 7.729579e-05, 5.720419e-07, -9.738964e-07, 2.1562724e-05, 7.707322e-05, 1.70712e-06, -9.141121e-07, -1.6732654e-05, 7.596262e-05, 2.802946e-06, -8.446863e-07, -5.425622e-05, 7.399141e-05, 3.8474677e-06, -7.6659353e-07, -9.058652e-05, 7.119654e-05, 4.82943e-06, -6.808917e-07, -0.00012532285, 6.762388e-05, 5.7384927e-06, -5.887091e-07, -0.0001580895, 6.332756e-05, 6.565335e-06, -4.912297e-07, -0.00018853977, 5.8369184e-05, 7.3017445e-06, -3.8967877e-07, -0.00021635942, 5.2817e-05, 7.940697e-06, -2.8530778e-07, -0.00024126982, 4.6744997e-05, 8.476415e-06, -1.7937968e-07, -0.00026303058, 4.0231964e-05, 8.904414e-06, -7.3153934e-08, -0.00028144172, 3.3360477e-05, 9.221534e-06, 3.2127932e-08, -0.00029634527, 2.6215896e-05, 9.425953e-06, 1.3525641e-07, -0.00030762635, 1.8885325e-05, 9.517186e-06, 2.350675e-07, -0.00031521395, 1.1456575e-05, 9.496067e-06, 3.3045538e-07, -0.0003190809, 4.017131e-06, 9.3647195e-06, 4.2038428e-07, -0.00031924344, -3.3468475e-06, 9.126507e-06, 5.038993e-07, -0.00031576038, -1.0551507e-05, 8.785978e-06, 5.80136e-07, -0.00030873172, -1.7516233e-05, 8.348788e-06, 6.48329e-07, -0.00029829674, -2.4164523e-05, 7.821619e-06, 7.0781925e-07, -0.00028463174, -3.042481e-05, 7.2120833e-06, 7.580597e-07, -0.00026794747, -3.6231206e-05, 6.5286226e-06, 7.9861974e-07, -0.00024848603, -4.152417e-05, 5.7803913e-06, 8.291885e-07, -0.0002265176, -4.625109e-05, 4.9771434e-06, 8.4957605e-07, -0.0002023368, -5.036678e-05, 4.1291064e-06, 8.597141e-07, -0.00017625892, -5.383387e-05, 3.2468565e-06, 8.59654e-07, -0.00014861595, -5.6623125e-05, 2.3411897e-06, 8.4956497e-07, -0.00011975233, -5.8713624e-05, 1.4229928e-06, 8.2972946e-07, -9.002095e-05, -6.0092883e-05, 5.031167e-07, 8.005384e-07, -5.977878e-05, -6.0756858e-05, -4.0774938e-07, 7.624847e-07, -2.9382736e-05, -6.0709834e-05, -1.2991989e-06, 7.161559e-07, 8.14462e-07, -5.9964248e-05, -2.1612236e-06, 6.622257e-07, 3.0468289e-05, -5.8540416e-05, -2.9843227e-06, 6.0144475e-07, 5.9246275e-05, -5.6466146e-05, -3.7596046e-06, 5.346306e-07, 8.6831635e-05, -5.377632e-05, -4.4788794e-06, 4.6265728e-07, 0.000112926675, -5.0512335e-05, -5.1347433e-06, 3.86444e-07, 0.00013725593, -4.6721547e-05, -5.7206485e-06, 3.0694392e-07, 0.00015956897, -4.2456617e-05, -6.230967e-06, 2.2513252e-07, 0.00017964284, -3.777479e-05, -6.6610396e-06, 1.4199584e-07, 0.00019728423, -3.2737193e-05, -7.0072147e-06, 5.8518935e-08, 0.0002123312, -2.7408027e-05, -7.2668718e-06, -2.4325521e-08, 0.00022465452, -2.1853803e-05, -7.438435e-06, -1.0558829e-07, 0.00023415861, -1.6142507e-05, -7.5213766e-06, -1.8435419e-07, 0.00024078209, -1.0342813e-05, -7.516201e-06, -2.597521e-07, 0.0002444979, -4.523257e-06, -7.4244263e-06, -3.3096438e-07, 0.0002453131, 1.2485418e-06, -7.2485464e-06, -3.9723534e-07, 0.00024326815, 6.9066514e-06, -6.991987e-06, -4.5787905e-07, 0.00023843585, 1.2387563e-05, -6.6590515e-06, -5.1228614e-07, 0.00023092006, 1.7630884e-05, -6.2548543e-06, -5.599294e-07, 0.0002208539, 2.2579985e-05, -5.7852503e-06, -6.0036876e-07, 0.00020839775, 2.718259e-05, -5.256753e-06, -6.3325484e-07, 0.0001937369, 3.139131e-05, -4.676449e-06, -6.583313e-07, 0.00017707904, 3.516412e-05, -4.051906e-06, -6.754366e-07, 0.00015865147, 3.846473e-05, -3.3910783e-06, -6.84504e-07, 0.00013869806, 4.1262923e-05, -2.702206e-06, -6.8556096e-07, 0.00011747629, 4.3534823e-05, -1.9937172e-06, -6.78727e-07, 9.5253905e-05, 4.526303e-05, -1.274126e-06, -6.642111e-07, 7.2305746e-05, 4.6436733e-05, -5.5193306e-07, -6.423075e-07, 4.891038e-05, 4.705172e-05, 1.6447315e-07, -6.133911e-07, 2.5346864e-05, 4.7110312e-05, 8.6691074e-07, -5.779116e-07, 1.8914722e-06, 4.662124e-05, 1.5474963e-06, -5.363872e-07, -2.1185442e-05, 4.559942e-05, 2.1987307e-06, -4.893973e-07, -4.3622476e-05, 4.4065688e-05, 2.81358e-06, -4.375749e-07, -6.517005e-05, 4.204645e-05, 3.3855483e-06, -3.815984e-07, -8.55931e-05, 3.9573297e-05, 3.9087445e-06, -3.2218284e-07, -0.00010467357, 3.668254e-05, 4.37794e-06, -2.6007118e-07, -0.00012221262, 3.341471e-05, 4.788619e-06, -1.9602507e-07, -0.00013803263, 2.9814035e-05, 5.137018e-06, -1.3081595e-07, -0.00015197888, 2.5927835e-05, 5.420156e-06, -6.521575e-08, -0.000163921, 2.1805956e-05, 5.6358576e-06, 1.1952672e-11, -0.000173754, 1.7500131e-05, 5.7827638e-06, 6.4120634e-08, -0.00018139913, 1.3063353e-05, 5.860334e-06, 1.263892e-07, -0.0001868043, 8.549245e-06, 5.8688393e-06, 1.8612985e-07, -0.00018994427, 4.011421e-06, 5.8093447e-06, 2.4269556e-07, -0.00019082046, -4.971275e-07, 5.683684e-06, 2.9548684e-07, -0.00018946052, -4.924638e-06, 5.494426e-06, 3.4395785e-07, -0.00018591754, -9.221154e-06, 5.2448327e-06, 3.8762184e-07, -0.00018026902, -1.3339076e-05, 4.9388077e-06, 4.2605583e-07, -0.0001726156, -1.7233668e-05, 4.580844e-06, 4.589044e-07, -0.00016307941, -2.0863534e-05, 4.1759586e-06, 4.8588265e-07, -0.00015180242, -2.4191033e-05, 3.7296281e-06, 5.0677835e-07, -0.00013894434, -2.7182663e-05, 3.2477167e-06, 5.214532e-07, -0.00012468056, -2.9809366e-05, 2.7364015e-06, 5.2984313e-07, -0.00010919985, -3.2046803e-05, 2.202096e-06, 5.319579e-07, -9.27019e-05, -3.3875545e-05, 1.651373e-06, 5.278795e-07, -7.5394855e-05, -3.5281228e-05, 1.090884e-06, 5.177603e-07, -5.7492776e-05, -3.625462e-05, 5.272819e-07, 5.018201e-07, -3.921303e-05, -3.679166e-05, -3.285569e-08, 4.803421e-07, -2.0773752e-05, -3.6893394e-05, -5.83102e-07, 4.5366892e-07, -2.3912733e-06, -3.6565907e-05, -1.1172526e-06, 4.221975e-07, 1.5722333e-05, -3.5820143e-05, -1.6293935e-06, 3.8637359e-07, 3.336164e-05, -3.4671713e-05, -2.113965e-06, 3.466858e-07, 5.033014e-05, -3.3140623e-05, -2.5658196e-06, 3.0365925e-07, 6.644237e-05, -3.1250976e-05, -2.9802754e-06, 2.5784885e-07, 8.152586e-05, -2.9030636e-05, -3.3531614e-06, 2.0983232e-07, 9.542295e-05, -2.6510814e-05, -3.6808583e-06, 1.6020327e-07, 0.00010799231, -2.3725677e-05, -3.960331e-06, 1.0956389e-07, 0.00011911037, -2.0711894e-05, -4.189153e-06, 5.8517998e-08, 0.0001286724, -1.750816e-05, -4.365525e-06, 7.663899e-09, 0.00013659344, -1.41547325e-05, -4.488286e-06, -4.2412374e-08, 0.00014280893, -1.0692924e-05, -4.556914e-06, -9.114367e-08, 0.00014727515, -7.1646145e-06, -4.5715233e-06, -1.3798794e-07, 0.00014996933, -3.6117533e-06, -4.5328516e-06, -1.8243412e-07, 0.00015088962, -7.587294e-08, -4.4422413e-06, -2.2400754e-07, 0.00015005471, 3.4023838e-06, -4.301613e-06, -2.622747e-07, 0.0001475033, 6.7837195e-06, -4.1134344e-06, -2.968478e-07, 0.00014329332, 1.0030616e-05, -3.880684e-06, -3.2738822e-07, 0.00013750092, 1.3107738e-05, -3.6068036e-06, -3.536098e-07, 0.00013021928, 1.5982303e-05, -3.2956561e-06, -3.752812e-07, 0.00012155731, 1.8624423e-05, -2.9514704e-06, -3.9222766e-07, 0.00011163802, 2.1007401e-05, -2.5787865e-06, -4.043321e-07, 0.00010059696, 2.3107985e-05, -2.182399e-06, -4.1153544e-07, 8.8580375e-05, 2.4906572e-05, -1.7672962e-06, -4.138364e-07, 7.574336e-05, 2.6387395e-05, -1.3386002e-06, -4.1129053e-07, 6.2247935e-05, 2.7538621e-05, -9.0150434e-07, -4.0400852e-07, 4.826102e-05, 2.8352426e-05, -4.6121215e-07, -3.9215408e-07, 3.395243e-05, 2.8825028e-05, -2.2877371e-08, -3.759412e-07, 1.9492882e-05, 2.8956656e-05, 4.0845538e-07, -3.5563068e-07, 5.0519816e-06, 2.8751478e-05, 8.279069e-07, -3.315265e-07, -9.203712e-06, 2.8217493e-05, 1.2308172e-06, -3.0397143e-07, -2.3112565e-05, 2.7366372e-05, 1.6127958e-06, -2.7334247e-07, -3.6519654e-05, 2.6213258e-05, 1.9697682e-06, -2.4004595e-07, -4.9278453e-05, 2.4776538e-05, 2.298017e-06, -2.045123e-07, -6.125238e-05, 2.3077575e-05, 2.5942204e-06, -1.6719062e-07, -7.2316216e-05, 2.1140404e-05, 2.8554823e-06, -1.2854323e-07, -8.2357365e-05, 1.8991419e-05, 3.0793606e-06, -8.904007e-08, -9.127695e-05, 1.6659023e-05, 3.2638857e-06, -4.9153147e-08, -9.899071e-05, 1.4173269e-05, 3.4075777e-06, -9.350997e-09, -0.00010542977, 1.1565476e-05, 3.509453e-06, 2.9906634e-08, -0.000110541114, 8.8678535e-06, 3.5690296e-06, 6.8173996e-08, -0.000114288, 6.113115e-06, 3.5863227e-06, 1.05024256e-07, -0.00011665008, 3.3340827e-06, 3.561837e-06, 1.4005413e-07, -0.00011762337, 5.6331345e-07, 3.4965524e-06, 1.7288812e-07, -0.000117220006, -2.1672777e-06, 3.3919043e-06, 2.0318245e-07, -0.00011546787, -4.826775e-06, 3.2497605e-06, 2.306285e-07, -0.00011240995, -7.3856017e-06, 3.0723913e-06, 2.5495575e-07, -0.00010810364, -9.815843e-06, 2.8624365e-06, 2.7593435e-07, -0.00010261982, -1.2091539e-05, 2.6228697e-06, 2.9337704e-07, -9.604178e-05, -1.4188953e-05, 2.3569569e-06, 3.071406e-07, -8.8464105e-05, -1.608681e-05, 2.0682148e-06, 3.1712682e-07, -7.9991325e-05, -1.7766497e-05, 1.7603655e-06, 3.2328285e-07, -7.07366e-05, -1.9212242e-05, 1.4372904e-06, 3.256011e-07, -6.0820214e-05, -2.0411244e-05, 1.1029816e-06, 3.2411845e-07, -5.0368115e-05, -2.1353771e-05, 7.6149513e-07, 3.1891526e-07, -3.951032e-05, -2.203322e-05, 4.1690186e-07, 3.1011356e-07, -2.8379354e-05, -2.244615e-05, 7.3240784e-08, 2.97875e-07, -1.7108689e-05, -2.2592254e-05, -2.6552746e-07, 2.8239836e-07, -5.8311625e-06, -2.2474325e-05, -5.955651e-07, 2.6391652e-07, 5.322533e-06, -2.209816e-05, -9.131995e-07, 2.426933e-07, 1.6225336e-05, -2.1472451e-05, -1.2149629e-06, 2.1901977e-07, 2.6755224e-05, -2.0608632e-05, -1.4976296e-06, 1.9321064e-07, 3.6796537e-05, -1.95207e-05, -1.7582483e-06, 1.6559994e-07, 4.6241214e-05, -1.8225011e-05, -1.9941729e-06, 1.3653707e-07, 5.4989916e-05, -1.6740056e-05, -2.2030865e-06, 1.0638233e-07, 6.295303e-05, -1.5086201e-05, -2.3830241e-06, 7.550269e-08, 7.0051545e-05, -1.32854275e-05, -2.532389e-06, 4.4267367e-08, 7.621777e-05, -1.1361051e-05, -2.649965e-06, 1.3043507e-08, 8.139596e-05, -9.337426e-06, -2.7349233e-06, -1.7807992e-08, 8.554275e-05, -7.2396447e-06, -2.786828e-06, -4.7936574e-08, 8.862743e-05, -5.0932417e-06, -2.8056313e-06, -7.7005915e-08, 9.063209e-05, -2.9238838e-06, -2.7916708e-06, -1.04697556e-07, 9.1551665e-05, -7.5707374e-07, -2.7456565e-06, -1.3071431e-07, 9.1393704e-05, 1.3821424e-06, -2.6686582e-06, -1.5478335e-07, 9.017812e-05, 3.4694579e-06, -2.5620861e-06, -1.7665892e-07, 8.793673e-05, 5.481574e-06, -2.4276687e-06, -1.9612479e-07, 8.47127e-05, 7.396453e-06, -2.2674285e-06, -2.129962e-07, 8.055987e-05, 9.193553e-06, -2.0836526e-06, -2.271215e-07, 7.5541895e-05, 1.0854037e-05, -1.8788618e-06, -2.3838341e-07, 6.97314e-05, 1.2360969e-05, -1.6557786e-06, -2.4669964e-07, 6.320899e-05, 1.3699472e-05, -1.4172914e-06, -2.5202348e-07, 5.6062112e-05, 1.4856868e-05, -1.1664183e-06, -2.5434352e-07, 4.8384034e-05, 1.5822789e-05, -9.0627026e-07, -2.5368337e-07, 4.0272582e-05, 1.6589256e-05, -6.400135e-07, -2.501007e-07, 3.1828968e-05, 1.7150733e-05, -3.7083197e-07, -2.4368606e-07, 2.3156555e-05, 1.7504153e-05, -1.01890066e-07, -2.3456117e-07, 1.435963e-05, 1.7648905e-05, 1.6370362e-07, -2.2287718e-07, 5.5421697e-06, 1.7586804e-05, 4.229313e-07, -2.0881225e-07, -3.1933469e-06, 1.7322034e-05, 6.728994e-07, -1.9256915e-07, -1.1747107e-05, 1.686105e-05, 9.108701e-07, -1.743724e-07, -2.0023072e-05, 1.621247e-05, 1.1342902e-06, -1.5446543e-07, -2.7930024e-05, 1.5386946e-05, 1.3408177e-06, -1.3310733e-07, -3.5382545e-05, 1.4396995e-05, 1.5283455e-06, -1.1056968e-07, -4.2301916e-05, 1.32568275e-05, 1.6950215e-06, -8.7133124e-08, -4.861689e-05, 1.1982159e-05, 1.8392662e-06, -6.3084016e-08, -5.4264423e-05, 1.0589995e-05, 1.9597862e-06, -3.8711e-08, -5.9190246e-05, 9.0984195e-06, 2.0555842e-06, -1.430163e-08, -6.334936e-05, 7.5263633e-06, 2.1259661e-06, 9.860944e-09, -6.670639e-05, 5.893373e-06, 2.170543e-06, 3.350118e-08, -6.923584e-05, 4.219372e-06, 2.189232e-06, 5.6354196e-08, -7.092221e-05, 2.5244262e-06, 2.1822507e-06, 7.816867e-08, -7.176004e-05, 8.285087e-07, 2.1501103e-06, 9.8709506e-08, -7.175378e-05, -8.4873153e-07, 2.093605e-06, 1.1776031e-07, -7.091756e-05, -2.48819e-06, 2.0137973e-06, 1.3512555e-07, -6.92749e-05, -4.071519e-06, 1.9120018e-06, 1.5063247e-07, -6.685826e-05, -5.5813275e-06, 1.7897659e-06, 1.6413277e-07, -6.370851e-05, -7.0013675e-06, 1.648847e-06, 1.7550381e-07, -5.987432e-05, -8.316701e-06, 1.4911902e-06, 1.8464969e-07, -5.541149e-05, -9.513851e-06, 1.318901e-06, 1.9150185e-07, -5.038214e-05, -1.0580937e-05, 1.1342196e-06, 1.9601949e-07, -4.485392e-05, -1.150778e-05, 9.3949166e-07, 1.9818941e-07, -3.8899136e-05, -1.22859965e-05, 7.371402e-07, 1.9802593e-07, -3.2593794e-05, -1.2909061e-05, 5.296358e-07, 1.9557007e-07, -2.6016718e-05, -1.3372358e-05, 3.1946735e-07, 1.9088873e-07, -1.9248537e-05, -1.3673193e-05, 1.09112754e-07, 1.8407341e-07, -1.2370756e-05, -1.3810802e-05, -9.898927e-08, 1.7523885e-07, -5.4647835e-06, -1.3786319e-05, -3.0246696e-07, 1.645212e-07, 1.3890079e-06, -1.3602737e-05, -4.9904185e-07, 1.5207614e-07, 8.1121925e-06, -1.3264842e-05, -6.8655345e-07, 1.3807673e-07, 1.4629167e-05, -1.2779124e-05, -8.6298246e-07, 1.2271113e-07, 2.086798e-05, -1.2153676e-05, -1.0264716e-06, 1.0618019e-07, 2.67611e-05, -1.1398073e-05, -1.1753446e-06, 8.869485e-08, 3.2246127e-05, -1.05232375e-05, -1.3081221e-06, 7.047359e-08, 3.726643e-05, -9.541287e-06, -1.4235364e-06, 5.1739743e-08, 4.1771702e-05, -8.4653775e-06, -1.5205416e-06, 3.2718837e-08, 4.5718432e-05, -7.309533e-06, -1.5983226e-06, 1.36359475e-08, 4.907031e-05, -6.0884668e-06, -1.6563004e-06, -5.286898e-09, 5.1798514e-05, -4.8174015e-06, -1.6941349e-06, -2.3833246e-08, 5.388192e-05, -3.511883e-06, -1.711725e-06, -4.1794628e-08, 5.530722e-05, -2.1875971e-06, -1.7092055e-06, -5.8972827e-08, 5.606895e-05, -8.601836e-07, -1.6869421e-06, -7.518202e-08, 5.616941e-05, 4.5494357e-07, -1.6455224e-06, -9.0250715e-08, 5.561852e-05, 1.7427701e-06, -1.5857463e-06, -1.04023485e-07, 5.4433567e-05, 2.9888492e-06, -1.5086126e-06, -1.16362514e-07, 5.2638887e-05, 4.179459e-06, -1.4153046e-06, -1.2714888e-07, 5.026547e-05, 5.3017493e-06, -1.3071726e-06, -1.3628365e-07, 4.735048e-05, 6.343876e-06, -1.1857163e-06, -1.4368864e-07, 4.393673e-05, 7.29512e-06, -1.0525642e-06, -1.49307e-07, 4.0072082e-05, 8.145996e-06, -9.094535e-07, -1.5310354e-07, 3.580882e-05, 8.888336e-06, -7.582069e-07, -1.5506474e-07, 3.1202966e-05, 9.515367e-06, -6.0071125e-07, -1.5519853e-07, 2.6313564e-05, 1.0021764e-05, -4.3889403e-07, -1.535339e-07, 2.1201959e-05, 1.0403686e-05, -2.7470048e-07, -1.5012013e-07, 1.5931031e-05, 1.0658799e-05, -1.100708e-07, -1.4502596e-07, 1.0564455e-05, 1.0786274e-05, 5.3082175e-08, -1.3833844e-07, 5.1659445e-06, 1.07867745e-05, 2.1289476e-07, -1.3016155e-07, -2.0148215e-07, 1.0662422e-05, 3.675731e-07, -1.2061484e-07, -5.4762245e-06, 1.0416747e-05, 5.1541275e-07, -1.0983168e-07, -1.0598786e-05, 1.0054626e-05, 6.548171e-07, -9.795754e-08, -1.5512429e-05, 9.5822015e-06, 7.843136e-07, -8.514806e-08, -2.0163783e-05, 9.00679e-06, 9.025693e-07, -7.156713e-08, -2.450341e-05, 8.336776e-06, 1.0084035e-06, -5.7384813e-08, -2.8486307e-05, 7.5815014e-06, 1.1007993e-06, -4.2775305e-08, -3.2072356e-05, 6.7511364e-06, 1.1789118e-06, -2.7914819e-08, -3.5226698e-05, 5.8565506e-06, 1.2420762e-06, -1.29795295e-08, -3.7920065e-05, 4.9091745e-06, 1.2898115e-06, 1.8564684e-09, -4.012901e-05, 3.9208594e-06, 1.3218233e-06, 1.6423142e-08, -4.1836083e-05, 2.9037305e-06, 1.3380044e-06, 3.0556418e-08, -4.302994e-05, 1.8700448e-06, 1.3384324e-06, 4.4099988e-08, -4.370537e-05, 8.320446e-07, 1.3233658e-06, 5.6906977e-08, -4.386325e-05, -1.9818224e-07, 1.2932386e-06, 6.8841494e-08, -4.3510423e-05, -1.2088404e-06, 1.2486513e-06, 7.978004e-08, -4.265954e-05, -2.1885587e-06, 1.1903622e-06, 8.961266e-08, -4.1328803e-05, -3.1265147e-06, 1.1192752e-06, 9.82441e-08, -3.954166e-05, -4.01255e-06, 1.0364272e-06, 1.0559456e-07, -3.7326456e-05, -4.837278e-06, 9.42974e-07, 1.1160041e-07, -3.471601e-05, -5.5921782e-06, 8.4017483e-07, 1.1621466e-07, -3.1747168e-05, -6.269682e-06, 7.293758e-07, 1.1940719e-07, -2.8460314e-05, -6.863243e-06, 6.1199336e-07, 1.2116487e-07, -2.4898829e-05, -7.367396e-06, 4.8949624e-07, 1.2149137e-07, -2.1108548e-05, -7.777802e-06, 3.633879e-07, 1.2040688e-07, -1.713719e-05, -8.0912805e-06, 2.3518831e-07, 1.17947565e-07, -1.3033769e-05, -8.305825e-06, 1.0641632e-07, 1.14164905e-07, -8.848008e-06, -8.42061e-06, -2.1428088e-08, 1.0912485e-07, -4.6297487e-06, -8.435976e-06, -1.4688077e-07, 1.02906775e-07, -4.283758e-07, -8.353412e-06, -2.6852976e-07, 9.5602374e-08, 3.7077489e-06, -8.1755115e-06, -3.8503077e-07, 8.731437e-08, 7.731828e-06, -7.905931e-06, -4.9512164e-07, 7.815517e-08, 1.1599147e-05, -7.5493263e-06, -5.9763545e-07, 6.824535e-08, 1.5267551e-05, -7.1112827e-06, -6.9151264e-07, 5.7712192e-08, 1.8697896e-05, -6.5982344e-06, -7.758113e-07, 4.668803e-08, 2.1854452e-05, -6.0173766e-06, -8.497161e-07, 3.5308684e-08, 2.4705249e-05, -5.3765684e-06, -9.125458e-07, 2.3711806e-08, 2.7222399e-05, -4.6842315e-06, -9.637586e-07, 1.2035253e-08, 2.938234e-05, -3.949244e-06, -1.0029563e-06, 4.1550688e-10, 3.1166037e-05, -3.1808268e-06, -1.0298866e-06, -1.10139e-08, 3.255914e-05, -2.3884359e-06, -1.0444431e-06, -2.2123873e-08, 3.3552045e-05, -1.5816453e-06, -1.0466648e-06, -3.2791178e-08, 3.4139954e-05, -7.7003534e-07, -1.0367326e-06, -4.2899764e-08, 3.432283e-05, 3.69178e-08, -1.0149648e-06, -5.2341996e-08, 3.410533e-05, 8.2995075e-07, -9.818118e-07, -6.1019755e-08, 3.349667e-05, 1.6001162e-06, -9.378482e-07, -6.88454e-08, 3.251043e-05, 2.3388816e-06, -8.8376385e-07, -7.574265e-08, 3.1164345e-05, 3.03822e-06, -8.2035433e-07, -8.1647215e-08, 2.948001e-05, 3.6906963e-06, -7.485099e-07, -8.650739e-08, 2.7482578e-05, 4.2895413e-06, -6.692034e-07, -9.028442e-08, 2.5200407e-05, 4.82872e-06, -5.83478e-07, -9.295275e-08, 2.2664673e-05, 5.3029903e-06, -4.9243346e-07, -9.450006e-08, 1.9908968e-05, 5.707948e-06, -3.972128e-07, -9.492723e-08, 1.696887e-05, 6.0400644e-06, -2.9898823e-07, -9.424809e-08, 1.3881489e-05, 6.2967147e-06, -1.989471e-07, -9.248904e-08, 1.0685027e-05, 6.4761903e-06, -9.827793e-08, -8.968854e-08, 7.4183044e-06, 6.5777053e-06, 1.8434313e-09, -8.589646e-08, 4.120308e-06, 6.6013895e-06, 1.0026714e-07, -8.117331e-08, 8.2973276e-07, 6.54827e-06, 1.9588225e-07, -7.558938e-08, -2.4154588e-06, 6.4202472e-06, 2.8762895e-07, -6.9223724e-08, -5.5784653e-06, 6.220056e-06, 3.7450994e-07, -6.216313e-08, -8.624052e-06, 5.951222e-06, 4.5560094e-07, -5.4500983e-08, -1.1518933e-05, 5.618005e-06, 5.3006016e-07, -4.6336062e-08, -1.4232124e-05, 5.225339e-06, 5.971367e-07, -3.777131e-08, -1.6735263e-05, 4.7787644e-06, 6.5617763e-07, -2.8912583e-08, -1.900289e-05, 4.2843517e-06, 7.0663407e-07, -1.9867352e-08, -2.1012702e-05, 3.7486245e-06, 7.4806553e-07, -1.0743461e-08, -2.2745751e-05, 3.178475e-06, 7.801436e-07, -1.6478545e-09, -2.4186611e-05, 2.5810787e-06, 8.026534e-07, 7.314643e-09, -2.5323492e-05, 1.9638057e-06, 8.1549456e-07, 1.6042502e-08, -2.6148327e-05, 1.334134e-06, 8.186803e-07, 2.4438608e-08, -2.6656788e-05, 6.99559e-07, 8.1233526e-07, 3.2411315e-08, -2.6848285e-05, 6.750777e-08, 7.966925e-07, 3.987541e-08, -2.672591e-05, -5.5474624e-07, 7.7208864e-07, 4.6752994e-08, -2.629633e-05, -1.1601646e-06, 7.3895853e-07, 5.297427e-08, -2.5569658e-05, -1.7420219e-06, 6.9782834e-07, 5.8478193e-08, -2.4559278e-05, -2.2939776e-06, 6.493081e-07, 6.321305e-08, -2.3281635e-05, -2.8101433e-06, 5.940831e-07, 6.713691e-08, -2.1755988e-05, -3.2851442e-06, 5.3290483e-07, 7.021791e-08, -2.0004149e-05, -3.7141713e-06, 4.665811e-07, 7.243448e-08, -1.8050176e-05, -4.093028e-06, 3.9596574e-07, 7.377544e-08, -1.5920072e-05, -4.4181697e-06, 3.21948e-07, 7.42399e-08, -1.3641439e-05, -4.686732e-06, 2.454416e-07, 7.3837164e-08, -1.1243135e-05, -4.8965535e-06, 1.6737378e-07, 7.2586396e-08, -8.754923e-06, -5.046189e-06, 8.8674355e-08, 7.0516265e-08, -6.2071076e-06, -5.134914e-06, 1.0264847e-08, 6.766444e-08, -3.630174e-06, -5.162721e-06, -6.6951976e-08, 6.407701e-08, -1.0544359e-06, -5.1303095e-06, -1.4210227e-07, 5.980781e-08, 1.4903147e-06, -5.0390613e-06, -2.1435072e-07, 5.4917674e-08, 3.9751435e-06, -4.8910183e-06, -2.829096e-07, 4.947358e-08, 6.3722937e-06, -4.6888445e-06, -3.4704712e-07, 4.354783e-08, 8.655489e-06, -4.435787e-06, -4.060948e-07, 3.721706e-08, 1.08002105e-05, -4.1356266e-06, -4.594544e-07, 3.056134e-08, 1.2783956e-05, -3.792626e-06, -5.0660344e-07, 2.3663135e-08, 1.4586458e-05, -3.411473e-06, -5.471001e-07, 1.660636e-08, 1.6189892e-05, -2.9972182e-06, -5.8058697e-07, 9.475348e-09, 1.757903e-05, -2.5552106e-06, -6.067938e-07, 2.3538813e-09, 1.8741386e-05, -2.091031e-06, -6.2553903e-07, -4.675767e-09, 1.9667305e-05, -1.6104239e-06, -6.3673053e-07, -1.1533766e-08, 2.0350028e-05, -1.1192269e-06, -6.403653e-07, -1.8143606e-08, 2.0785727e-05, -6.233033e-07, -6.365276e-07, -2.4432934e-08, 2.0973497e-05, -1.2847242e-07, -6.2538703e-07, -3.0334313e-08, 2.0915319e-05, 3.5955634e-07, -6.071947e-07, -3.5785927e-08, 2.0615984e-05, 8.3524793e-07, -5.8227926e-07, -4.0732203e-08, 2.0082998e-05, 1.2933027e-06, -5.510416e-07, -4.512434e-08, 1.9326444e-05, 1.7287141e-06, -5.139491e-07, -4.8920786e-08, 1.8358827e-05, 2.136821e-06, -4.7152912e-07, -5.208755e-08, 1.719488e-05, 2.513357e-06, -4.2436182e-07, -5.459853e-08, 1.5851365e-05, 2.854492e-06, -3.730726e-07, -5.6435628e-08, 1.4346844e-05, 3.1568707e-06, -3.1832414e-07, -5.7588863e-08, 1.2701429e-05, 3.417641e-06, -2.6080804e-07, -5.805633e-08, 1.0936526e-05, 3.6344818e-06, -2.0123633e-07, -5.784409e-08, 9.074568e-06, 3.8056182e-06, -1.40333e-07, -5.6965984e-08, 7.138734e-06, 3.9298347e-06, -7.882523e-08, -5.544332e-08, 5.152669e-06, 4.0064797e-06, -1.7435102e-08, -5.33045e-08, 3.1402064e-06, 4.0354616e-06, 4.312879e-08, -5.0584603e-08, 1.1250844e-06, 4.0172436e-06, 1.02179264e-07, -4.7324832e-08, -8.693256e-07, 3.9528263e-06, 1.5905817e-07, -4.3571955e-08, -2.8202828e-06, 3.8437292e-06, 2.131435e-07, -3.937766e-08, -4.70593e-06, 3.6919637e-06, 2.6385598e-07, -3.4797885e-08, -6.5055324e-06, 3.5000005e-06, 3.1066514e-07, -2.9892096e-08, -8.199699e-06, 3.2707346e-06, 3.530945e-07, -2.4722523e-08, -9.770581e-06, 3.0074448e-06, 3.9072623e-07, -1.935342e-08, -1.120206e-05, 2.713748e-06, 4.2320514e-07, -1.3850275e-08, -1.2479897e-05, 2.3935534e-06, 4.5024154e-07, -8.279025e-09, -1.3591873e-05, 2.0510108e-06, 4.7161362e-07, -2.705293e-09, -1.4527891e-05, 1.6904595e-06, 4.8716885e-07, 2.8063643e-09, -1.5280062e-05, 1.3163748e-06, 4.9682455e-07, 8.193193e-09, -1.5842756e-05, 9.3331323e-07, 5.005677e-07, 1.3394932e-08, -1.6212629e-05, 5.4585934e-07, 4.984541e-07, 1.8354473e-08, -1.6388629e-05, 1.585717e-07, 4.906061e-07, 2.3018469e-08, -1.6371963e-05, -2.2406947e-07, 4.772107e-07, 2.7337883e-08, -1.6166048e-05, -5.9771264e-07, 4.5851576e-07, 3.1268492e-08, -1.5776437e-05, -9.581833e-07, 4.3482646e-07, 3.4771308e-08, -1.5210711e-05, -1.3015293e-06, 4.0650062e-07, 3.781295e-08, -1.447837e-05, -1.624063e-06, 3.7394372e-07, 4.036594e-08, -1.3590677e-05, -1.9223992e-06, 3.376035e-07, 4.2408903e-08, -1.2560508e-05, -2.1934895e-06, 2.9796394e-07, 4.392674e-08, -1.1402173e-05, -2.434652e-06, 2.5553908e-07, 4.4910674e-08, -1.0131225e-05, -2.6435964e-06, 2.1086669e-07, 4.5358256e-08, -8.76426e-06, -2.818443e-06, 1.6450147e-07, 4.527329e-08, -7.31871e-06, -2.9577386e-06, 1.1700846e-07, 4.4665676e-08, -5.8126207e-06, -3.060466e-06, 6.895629e-08, 4.35512e-08, -4.26444e-06, -3.1260481e-06, 2.0910543e-08, 4.195125e-08, -2.692793e-06, -3.1543477e-06, -2.6572744e-08, 3.9892477e-08, -1.1162645e-06, -3.1456611e-06, -7.295335e-08, 3.7406398e-08, 4.4681502e-07, -3.100708e-06, -1.17712865e-07, 3.452894e-08, 1.9785773e-06, -3.0206158e-06, -1.6036032e-07, 3.1299972e-08, 3.4618163e-06, -2.9068997e-06, -2.0043741e-07, 2.7762754e-08, 4.8801753e-06, -2.7614387e-06, -2.3752328e-07, 2.3963391e-08, 6.2183217e-06, -2.586448e-06, -2.712387e-07, 1.9950253e-08, 7.4621094e-06, -2.3844475e-06, -3.0124983e-07, 1.5773377e-08, 8.59872e-06, -2.1582275e-06, -3.2727132e-07, 1.148385e-08, 9.616792e-06, -1.9108118e-06, -3.4906873e-07, 7.133216e-09, 1.0506524e-05, -1.645419e-06, -3.6646045e-07, 2.772857e-09, 1.12597645e-05, -1.3654222e-06, -3.7931895e-07, -1.5465892e-09, 1.1870081e-05, -1.0743067e-06, -3.8757128e-07, -5.7758074e-09, 1.23328e-05, -7.756284e-07, -3.91199e-07, -9.867353e-09, 1.2645036e-05, -4.72971e-07, -3.9023757e-07, -1.3776168e-08, 1.2805693e-05, -1.6990451e-07, -3.8477492e-07, -1.7460064e-08, 1.2815448e-05, 1.3005625e-07, -3.7494965e-07, -2.0880165e-08, 1.2676715e-05, 4.234912e-07, -3.6094852e-07, -2.4001295e-08, 1.2393585e-05, 7.07113e-07, -3.4300348e-07, -2.6792332e-08, 1.19717515e-05, 9.77803e-07, -3.213883e-07, -2.9226493e-08, 1.1418419e-05, 1.2326444e-06, -2.9641464e-07, -3.1281576e-08, 1.0742192e-05, 1.4689527e-06, -2.6842778e-07, -3.294014e-08, 9.952956e-06, 1.6843028e-06, -2.3780213e-07, -3.418962e-08, 9.061738e-06, 1.8765529e-06, -2.0493634e-07, -3.5022403e-08, 8.0805585e-06, 2.0438645e-06, -1.7024837e-07, -3.543582e-08, 7.022283e-06, 2.1847181e-06, -1.3417024e-07, -3.5432116e-08, 5.90045e-06, 2.2979264e-06, -9.714284e-08, -3.5018306e-08, 4.7291087e-06, 2.382642e-06, -5.961066e-08, -3.420605e-08, 3.522645e-06, 2.4383608e-06, -2.201661e-08, -3.3011418e-08, 2.2956121e-06, 2.4649235e-06, 1.5203117e-08, -3.145464e-08, 1.0625567e-06, 2.4625108e-06, 5.1623957e-08, -2.95598e-08, -1.6214814e-07, 2.4316355e-06, 8.68377e-08, -2.7354488e-08, -1.3644666e-06, 2.3731318e-06, 1.2045693e-07, -2.486943e-08, -2.5308568e-06, 2.2881388e-06, 1.5211921e-07, -2.2138071e-08, -3.6484198e-06, 2.1780843e-06, 1.8149078e-07, -1.9196154e-08, -4.7050376e-06, 2.0446614e-06, 2.0827e-07, -1.6081255e-08, -5.6894996e-06, 1.8898058e-06, 2.3219027e-07, -1.2832329e-08, -6.59162e-06, 1.7156688e-06, 2.530226e-07, -9.489224e-09, -7.402335e-06, 1.5245887e-06, 2.7057752e-07, -6.0922143e-09, -8.113791e-06, 1.319061e-06, 2.847067e-07, -2.6815246e-09, -8.719416e-06, 1.1017064e-06, 2.953039e-07, 7.031364e-10, -9.21397e-06, 8.75239e-07, 3.0230558e-07, 4.023026e-09, -9.593588e-06, 6.4243255e-07, 3.0569092e-07, 7.240799e-09, -9.855804e-06, 4.0608802e-07, 3.0548125e-07, 1.0320919e-08, -9.999545e-06, 1.6900032e-07, 3.0173916e-07, 1.3230036e-08, -1.0025133e-05, -6.6073824e-08, 2.945671e-07, 1.5937339e-08, -9.934248e-06, -2.964471e-07, 2.841055e-07, 1.8414866e-08, -9.729894e-06, -5.195316e-07, 2.7053053e-07, 2.0637788e-08, -9.416336e-06, -7.328672e-07, 2.5405143e-07, 2.2584635e-08, -8.999032e-06, -9.3414764e-07, 2.3490755e-07, 2.423749e-08, -8.484549e-06, -1.121245e-06, 2.1336508e-07, 2.5582146e-08, -7.88047e-06, -1.2922309e-06, 1.8971357e-07, 2.6608195e-08, -7.195287e-06, -1.445396e-06, 1.6426205e-07, 2.7309092e-08, -6.4382893e-06, -1.5792658e-06, 1.3733528e-07, 2.7682168e-08, -5.6194417e-06, -1.6926138e-06, 1.0926961e-07, 2.772859e-08, -4.7492586e-06, -1.7844712e-06, 8.040899e-08, 2.745329e-08, -3.8386715e-06, -1.854135e-06, 5.110077e-08, 2.6864837e-08, -2.8988977e-06, -1.9011702e-06, 2.16917e-08, 2.5975288e-08, -1.9413042e-06, -1.9254112e-06, -7.476121e-09, 2.4799975e-08, -9.772733e-07, -1.926959e-06, -3.6069117e-08, 2.335729e-08, -1.807226e-08, -1.9061755e-06, -6.3765945e-08, 2.1668402e-08, 9.252769e-07, -1.8636753e-06, -9.026101e-08, 1.9756987e-08, 1.8421199e-06, -1.800314e-06, -1.1526775e-07, 1.764889e-08, 2.7222877e-06, -1.717174e-06, -1.3852163e-07, 1.5371805e-08, 3.5562061e-06, -1.6155491e-06, -1.5978283e-07, 1.295492e-08, 4.3349964e-06, -1.4969248e-06, -1.788386e-07, 1.0428548e-08, 5.0505664e-06, -1.3629591e-06, -1.9550531e-07, 7.823766e-09, 5.695692e-06, -1.2154594e-06, -2.0963e-07, 5.172035e-09, 6.264085e-06, -1.0563596e-06, -2.2109177e-07, 2.504836e-09, 6.75045e-06, -8.8769553e-07, -2.2980251e-07, -1.4670004e-10, 7.150531e-06, -7.115797e-07, -2.3570743e-07, -2.7521438e-09, 7.4611416e-06, -5.301753e-07, -2.387852e-07, -5.282109e-09, 7.680183e-06, -3.456709e-07, -2.3904747e-07, -7.708576e-09, 7.806654e-06, -1.6025395e-07, -2.3653838e-07, -1.000519e-08, 7.840639e-06, 2.391398e-08, -2.3133336e-07, -1.2147542e-08, 7.783295e-06, 2.0472201e-07, -2.2353777e-07, -1.4113417e-08, 7.636812e-06, 3.8013349e-07, -2.1328523e-07, -1.5883016e-08, 7.40438e-06, 5.482083e-07, -2.0073556e-07, -1.7439138e-08, 7.090127e-06, 7.071237e-07, -1.8607247e-07, -1.876735e-08, 6.699061e-06, 8.5519366e-07, -1.6950105e-07, -1.985609e-08, 6.2369945e-06, 9.908856e-07, -1.5124509e-07, -2.0696767e-08, 5.7104644e-06, 1.1128363e-06, -1.315441e-07, -2.1283801e-08, 5.1266447e-06, 1.219864e-06, -1.1065032e-07, -2.1614644e-08, 4.4932526e-06, 1.3109797e-06, -8.882555e-08, -2.168976e-08, 3.8184494e-06, 1.385395e-06, -6.633802e-08, -2.1512554e-08, 3.1107395e-06, 1.4425282e-06, -4.3459114e-08, -2.1089306e-08, 2.3788657e-06, 1.4820073e-06, -2.046021e-08, -2.0429034e-08, 1.6317043e-06, 1.5036707e-06, 2.390464e-09, -1.9543348e-08, 8.781599e-07, 1.5075659e-06, 2.4830888e-08, -1.8446276e-08, 1.2706168e-07, 1.4939454e-06, 4.6608175e-08, -1.7154052e-08, -6.12937e-07, 1.4632601e-06, 6.748136e-08, -1.5684906e-08, -1.3334562e-06, 1.4161506e-06, 8.722395e-08, -1.4058801e-08, -2.0264818e-06, 1.3534374e-06, 1.0562636e-07, -1.229719e-08, -2.684452e-06, 1.2761074e-06, 1.2249802e-07, -1.0422732e-08, -3.3003373e-06, 1.1853006e-06, 1.3766926e-07, -8.459013e-09, -3.8677135e-06, 1.0822936e-06, 1.5099292e-07, -6.430259e-09, -4.3808245e-06, 9.68483e-07, 1.6234573e-07, -4.3610413e-09, -4.8346396e-06, 8.453671e-07, 1.7162925e-07, -2.2759892e-09, -5.2248984e-06, 7.145266e-07, 1.7877069e-07, -1.9950301e-10, -5.548147e-06, 5.776055e-07, 1.8372322e-07, 1.844525e-09, -5.801766e-06, 4.362903e-07, 1.8646618e-07, 3.832978e-09, -5.9839845e-06, 2.9229045e-07, 1.8700479e-07, 5.7437695e-09, -6.093889e-06, 1.4731768e-07, 1.8536974e-07, 7.556082e-09, -6.1314176e-06, 3.0663436e-09, 1.8161633e-07, 9.250585e-09, -6.097348e-06, -1.3880587e-07, 1.7582347e-07, 1.08096385e-08, -5.9932718e-06, -2.766966e-07, 1.6809237e-07, 1.2217463e-08, -5.8215664e-06, -4.090764e-07, 1.5854495e-07, 1.3460292e-08, -5.585351e-06, -5.3450515e-07, 1.4732214e-07, 1.4526505e-08, -5.28844e-06, -6.5164744e-07, 1.345819e-07, 1.5406716e-08, -4.935286e-06, -7.592859e-07, 1.2049708e-07, 1.6093848e-08, -4.5309184e-06, -8.563338e-07, 1.0525326e-07, 1.6583183e-08, -4.0808745e-06, -9.418451e-07, 8.904626e-08, 1.6872365e-08, -3.5911287e-06, -1.015023e-06, 7.2079835e-08, 1.69614e-08, -3.0680144e-06, -1.075227e-06, 5.4563067e-08, 1.6852606e-08, -2.518145e-06, -1.1219774e-06, 3.6707938e-08, 1.6550556e-08, -1.9483334e-06, -1.1549583e-06, 1.8726793e-08, 1.606198e-08, -1.3655091e-06, -1.1740184e-06, 8.2987467e-10, 1.5395658e-08, -7.766358e-07, -1.1791701e-06, -1.6777065e-08, 1.4562276e-08, -1.886312e-07, -1.1705865e-06, -3.3895077e-08, 1.3574279e-08, 3.9171306e-07, -1.1485972e-06, -5.0334197e-08, 1.2445691e-08, 9.578077e-07, -1.1136808e-06, -6.591551e-08, 1.1191929e-08, 1.5033388e-06, -1.066458e-06, -8.0473e-08, 9.829603e-09, 2.0223358e-06, -1.0076815e-06, -9.385532e-08, 8.376298e-09, 2.5092359e-06, -9.3822496e-07, -1.05927235e-07, 6.85036e-09, 2.95894e-06, -8.590712e-07, -1.1657094e-07, 5.270668e-09, 3.366866e-06, -7.712987e-07, -1.2568714e-07, 3.6564072e-09, 3.728991e-06, -6.760677e-07, -1.3319588e-07, 2.0268422e-09, 4.0418904e-06, -5.7460545e-07, -1.3903717e-07, 4.0109174e-10, 4.3027667e-06, -4.681907e-07, -1.4317129e-07, -1.2020895e-09, 4.5094707e-06, -3.581381e-07, -1.4557898e-07, -2.7645222e-09, 4.660517e-06, -2.457824e-07, -1.4626126e-07, -4.2688026e-09, 4.7550884e-06, -1.3246272e-07, -1.4523911e-07, -5.698492e-09, 4.7930366e-06, -1.9506862e-08, -1.4255292e-07, -7.0382895e-09, 4.7748695e-06, 9.178376e-08, -1.3826161e-07, -8.274192e-09, 4.7017375e-06, 2.0014883e-07, -1.3244174e-07, -9.393632e-09, 4.5754064e-06, 3.0438298e-07, -1.2518626e-07, -1.0385602e-08, 4.39823e-06, 4.0334885e-07, -1.1660318e-07, -1.1240753e-08, 4.17311e-06, 4.9598907e-07, -1.0681408e-07, -1.1951477e-08, 3.903455e-06, 5.8133725e-07, -9.595246e-08, -1.2511965e-08, 3.5931316e-06, 6.585275e-07, -8.4162e-08, -1.2918243e-08, 3.246413e-06, 7.268029e-07, -7.159472e-08, -1.3168191e-08, 2.8679215e-06, 7.8552245e-07, -5.8409096e-08, -1.3261532e-08, 2.4625701e-06, 8.3416637e-07, -4.4768104e-08, -1.3199808e-08, 2.0355008e-06, 8.723403e-07, -3.0837267e-08, -1.29863285e-08, 1.5920206e-06, 8.9977766e-07, -1.6782687e-08, -1.2626104e-08, 1.1375372e-06, 9.163406e-07, -2.7691178e-09, -1.2125762e-08, 6.7749596e-07, 9.220194e-07, 1.1041917e-08, -1.1493438e-08, 2.1731475e-07, 9.169306e-07, 2.4493941e-08, -1.0738662e-08, -2.3767731e-07, 9.0131334e-07, 3.7437257e-08, -9.872221e-09, -6.823005e-07, 8.755247e-07, 4.973056e-08, -8.906012e-09, -1.1115818e-06, 8.4003335e-07, 6.124243e-08, -7.852889e-09, -1.520809e-06, 7.954126e-07, 7.185271e-08, -6.7264976e-09, -1.9055809e-06, 7.423318e-07, 8.145366e-08, -5.5411027e-09, -2.2618533e-06, 6.8154696e-07, 8.995106e-08, -4.3114126e-09, -2.585979e-06, 6.1389073e-07, 9.726501e-08, -3.0524028e-09, -2.8747447e-06, 5.4026117e-07, 1.0333066e-07, -1.7791372e-09, -3.1253996e-06, 4.616106e-07, 1.0809872e-07, -5.065927e-10, -3.3356807e-06, 3.789335e-07, 1.115357e-07, 7.505129e-10, -3.5038295e-06, 2.9325426e-07, 1.13624104e-07, 1.9778867e-09, -3.628605e-06, 2.0561488e-07, 1.1436234e-07, 3.16182e-09, -3.709289e-06, 1.1706265e-07, 1.1376446e-07, 4.289335e-09, -3.745686e-06, 2.8637835e-08, 1.1185975e-07, 5.3483262e-09, -3.7381158e-06, -5.863815e-08, 1.08692134e-07, 6.3276815e-09, -3.687402e-06, -1.437743e-07, 1.0431943e-07, 7.2173987e-09, -3.5948542e-06, -2.2582097e-07, 9.8812414e-08, 8.00868e-09, -3.462244e-06, -3.0388017e-07, 9.225383e-08, 8.694013e-09, -3.2917767e-06, -3.771151e-07, 8.473719e-08, 9.267239e-09, -3.0860597e-06, -4.447588e-07, 7.6365545e-08, 9.723601e-09, -2.848064e-06, -5.061219e-07, 6.7250106e-08, 1.0059771e-08, -2.5810848e-06, -5.6059923e-07, 5.7508842e-08, 1.0273871e-08, -2.2886982e-06, -6.0767553e-07, 4.7264983e-08, 1.0365465e-08, -1.9747133e-06, -6.469297e-07, 3.664552e-08, 1.0335545e-08, -1.6431266e-06, -6.7803836e-07, 2.5779663e-08, 1.0186492e-08, -1.2980707e-06, -7.007778e-07, 1.479731e-08, 9.922023e-09, -9.4376543e-07, -7.1502484e-07, 3.827534e-09, 9.547135e-09, -5.8446665e-07, -7.2075676e-07, -7.002899e-09, 9.068013e-09, -2.2441691e-07, -7.180498e-07, -1.7570958e-08, 8.491949e-09, 1.3220347e-07, -7.0707654e-07, -2.7758706e-08, 7.827235e-09, 4.813239e-07, -6.8810243e-07, -3.7454587e-08, 7.0830475e-09, 8.190289e-07, -6.614809e-07, -4.65546e-08, 6.2693317e-09, 1.1416005e-06, -6.2764826e-07, -5.496339e-08, 5.3966707e-09, 1.445558e-06, -5.871168e-07, -6.25952e-08, 4.4761523e-09, 1.7276949e-06, -5.404678e-07, -6.937468e-08, 3.5192327e-09, 1.9851104e-06, -4.883437e-07, -7.5237644e-08, 2.537598e-09, 2.215239e-06, -4.3143942e-07, -8.013156e-08, 1.5430243e-09, 2.4158735e-06, -3.7049375e-07, -8.401601e-08, 5.472409e-10, 2.5851853e-06, -3.0627973e-07, -8.686292e-08, -4.3820567e-10, 2.7217388e-06, -2.395954e-07, -8.865671e-08, -1.4020818e-09, 2.824502e-06, -1.7125402e-07, -8.939425e-08, -2.3335915e-09, 2.8928507e-06, -1.02074345e-07, -8.908468e-08, -3.2224943e-09, 2.92657e-06, -3.2871213e-08, -8.774912e-08, -4.0592143e-09, 2.9258495e-06, 3.555395e-08, -8.54202e-08, -4.8349396e-09, 2.8912737e-06, 1.02422135e-07, -8.2141504e-08, -5.5417124e-09, 2.8238098e-06, 1.6698539e-07, -7.796689e-08, -6.172506e-09, 2.7247893e-06, 2.2853496e-07, -7.295968e-08, -6.7212906e-09, 2.5958864e-06, 2.8640886e-07, -6.719176e-08, -7.183087e-09, 2.4390934e-06, 3.3999873e-07, -6.074264e-08, -7.554006e-09, 2.2566924e-06, 3.8875592e-07, -5.3698376e-08, -7.831276e-09, 2.0512232e-06, 4.3219703e-07, -4.615046e-08, -8.013254e-09, 1.8254502e-06, 4.6990817e-07, -3.81947e-08, -8.0994305e-09, 1.582327e-06, 5.0154875e-07, -2.993001e-08, -8.09041e-09, 1.3249578e-06, 5.2685414e-07, -2.1457227e-08, -7.987892e-09, 1.0565604e-06, 5.456375e-07, -1.2877911e-08, -7.794628e-09, 7.804263e-07, 5.577906e-07, -4.2931516e-09, -7.514375e-09, 4.998811e-07, 5.6328366e-07, 4.1975903e-09, -7.151831e-09, 2.1824597e-07, 5.6216476e-07, 1.2497605e-08, -6.7125727e-09, -6.1200744e-08, 5.545574e-07, 2.0514012e-08, -6.2029675e-09, -3.352611e-07, 5.406583e-07, 2.8158766e-08, -5.630092e-09, -6.008529e-07, 5.207337e-07, 3.53496e-08, -5.0016364e-09, -8.5504377e-07, 4.9511505e-07, 4.201088e-08, -4.3258064e-09, -1.0950822e-06, 4.641942e-07, 4.807436e-08, -3.6112175e-09, -1.3184266e-06, 4.2841788e-07, 5.3479866e-08, -2.86679e-09, -1.5227712e-06, 3.8828145e-07, 5.817584e-08, -2.1016404e-09, -1.7060687e-06, 3.4432253e-07, 6.21198e-08, -1.3249726e-09, -1.8665498e-06, 2.971139e-07, 6.527869e-08, -5.459693e-10, -2.002739e-06, 2.4725642e-07, 6.762909e-08, 2.2631316e-10, -2.1134663e-06, 1.9537156e-07, 6.915731e-08, 9.83048e-10, -2.1978763e-06, 1.4209381e-07, 6.9859446e-08, 1.715736e-09, -2.2554327e-06, 8.806321e-08, 6.974118e-08, 2.4162987e-09, -2.2859185e-06, 3.391776e-08, 6.8817634e-08, 3.0771647e-09, -2.2894344e-06, -1.9713866e-08, 6.711297e-08, 3.6913492e-09, -2.266391e-06, -7.221948e-08, 6.465999e-08, 4.2525237e-09, -2.2174995e-06, -1.2301017e-07, 6.149963e-08, 4.7550803e-09, -2.1437586e-06, -1.7152672e-07, 5.76803e-08, 5.1941833e-09, -2.046438e-06, -2.1724563e-07, 5.3257242e-08, 5.565812e-09, -1.927059e-06, -2.5968453e-07, 4.8291767e-08, 5.8667937e-09, -1.7873724e-06, -2.9840706e-07, 4.2850427e-08, 6.0948278e-09, -1.6293353e-06, -3.3302726e-07, 3.7004174e-08, 6.248496e-09, -1.4550841e-06, -3.6321305e-07, 3.0827458e-08, 6.327264e-09, -1.2669072e-06, -3.8868924e-07, 2.4397309e-08, 6.331474e-09, -1.0672161e-06, -4.092398e-07, 1.7792399e-08, 6.2623253e-09, -8.585148e-07, -4.247093e-07, 1.1092104e-08, 6.121847e-09, -6.4336996e-07, -4.3500376e-07, 4.3755817e-09, 5.912858e-09, -4.2437983e-07, -4.4009064e-07, -2.2791529e-09, 5.6389258e-09, -2.0414359e-07, -4.3999825e-07, -8.796104e-09, 5.304307e-09, 1.47686166e-08, -4.3481432e-07, -1.5102144e-08, 4.913892e-09, 2.2984501e-07, -4.2468412e-07, -2.1127807e-08, 4.473133e-09, 4.3866027e-07, -4.098077e-07, -2.6808044e-08, 3.9879753e-09, 6.389021e-07, -3.9043675e-07, -3.208288e-08, 3.4647774e-09, 8.2839625e-07, -3.6687072e-07, -3.6898054e-08, 2.9102325e-09, 1.0051291e-06, -3.3945258e-07, -4.1205517e-08, 2.3312843e-09, 1.1672687e-06, -3.0856424e-07, -4.496391e-08, 1.7350429e-09, 1.3131826e-06, -2.7462127e-07, -4.8138922e-08, 1.128699e-09, 1.4414532e-06, -2.3806776e-07, -5.070357e-08, 5.194406e-10, 1.5508913e-06, -1.993705e-07, -5.2638377e-08, -8.563136e-11, 1.6405454e-06, -1.5901331e-07, -5.39315e-08, -6.795831e-10, 1.7097088e-06, -1.1749112e-07, -5.457871e-08, -1.2557257e-09, 1.7579241e-06, -7.530406e-08, -5.4583328e-08, -1.8076884e-09, 1.7849839e-06, -3.2951583e-08, -5.3956057e-08, -2.3294868e-09, 1.790929e-06, 9.073299e-09, -5.2714736e-08, -2.815586e-09, 1.7760442e-06, 5.028963e-08, -5.0884015e-08, -3.260957e-09, 1.7408503e-06, 9.023385e-08, -4.849495e-08, -3.6611263e-09, 1.686095e-06, 1.284649e-07, -4.5584542e-08, -4.0122186e-09, 1.6127392e-06, 1.6456893e-07, -4.2195207e-08, -4.3109916e-09, 1.5219435e-06, 1.9816363e-07, -3.8374196e-08, -4.5548623e-09};
endpackage
`endif
