`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam N = 4;
	localparam M = 4;
	localparam real Lfr[0:3] = {0.6944144, 0.6944144, 0.77749187, 0.77749187};
	localparam real Lfi[0:3] = {0.53008276, -0.53008276, 0.1975122, -0.1975122};
	localparam real Lbr[0:3] = {0.6944144, 0.6944144, 0.77749187, 0.77749187};
	localparam real Lbi[0:3] = {0.53008276, -0.53008276, 0.1975122, -0.1975122};
	localparam real Wfr[0:3] = {0.25414562, 0.25414562, -0.010946152, -0.010946152};
	localparam real Wfi[0:3] = {-0.019789157, 0.019789157, -0.25008067, 0.25008067};
	localparam real Wbr[0:3] = {-0.25414562, -0.25414562, -0.010946152, -0.010946152};
	localparam real Wbi[0:3] = {0.019789157, -0.019789157, -0.25008067, 0.25008067};
	localparam real Ffr[0:3][0:79] = '{
		'{0.17863393, -0.09251931, -0.25321913, 0.060769558, 0.094903484, -0.20938554, -0.12451469, 0.11594125, -0.0045285556, -0.22019, 0.020327035, 0.11464327, -0.07871964, -0.14600335, 0.12326026, 0.07073361, -0.10587191, -0.03472484, 0.15567382, 0.01074123, -0.08695919, 0.06320277, 0.12213215, -0.03906609, -0.039970078, 0.114279784, 0.050810527, -0.062453806, 0.010855579, 0.11047875, -0.022644024, -0.056922436, 0.045581665, 0.06621784, -0.07022722, -0.031390827, 0.05502016, 0.0076479567, -0.08025168, -0.00015333144, 0.041625693, -0.03991569, -0.05785849, 0.0237445, 0.015819622, -0.06127297, -0.019107524, 0.033094063, -0.009797943, -0.054634042, 0.017620465, 0.027840206, -0.025681186, -0.029113853, 0.039054655, 0.0134079205, -0.028188987, 0.0012624935, 0.0407923, -0.002626315, -0.019549819, 0.023973053, 0.026847044, -0.013880414, -0.00563754, 0.03233093, 0.0061533004, -0.017273117, 0.0070908256, 0.026605913, -0.011943759, -0.013395881, 0.014150508, 0.0122761205, -0.021284029, -0.005421758, 0.01424092, -0.0032561799, -0.020444404, 0.0026938305},
		'{0.17863393, -0.09251931, -0.25321913, 0.060769558, 0.094903484, -0.20938554, -0.12451469, 0.11594125, -0.0045285556, -0.22019, 0.020327035, 0.11464327, -0.07871964, -0.14600335, 0.12326026, 0.07073361, -0.10587191, -0.03472484, 0.15567382, 0.01074123, -0.08695919, 0.06320277, 0.12213215, -0.03906609, -0.039970078, 0.114279784, 0.050810527, -0.062453806, 0.010855579, 0.11047875, -0.022644024, -0.056922436, 0.045581665, 0.06621784, -0.07022722, -0.031390827, 0.05502016, 0.0076479567, -0.08025168, -0.00015333144, 0.041625693, -0.03991569, -0.05785849, 0.0237445, 0.015819622, -0.06127297, -0.019107524, 0.033094063, -0.009797943, -0.054634042, 0.017620465, 0.027840206, -0.025681186, -0.029113853, 0.039054655, 0.0134079205, -0.028188987, 0.0012624935, 0.0407923, -0.002626315, -0.019549819, 0.023973053, 0.026847044, -0.013880414, -0.00563754, 0.03233093, 0.0061533004, -0.017273117, 0.0070908256, 0.026605913, -0.011943759, -0.013395881, 0.014150508, 0.0122761205, -0.021284029, -0.005421758, 0.01424092, -0.0032561799, -0.020444404, 0.0026938305},
		'{-0.040811576, -0.16744499, -0.0013990296, -0.24659619, -0.08905777, -0.12068868, -0.035101686, -0.18322004, -0.11222095, -0.0799173, -0.053682268, -0.12621841, -0.117192656, -0.046606373, -0.060886957, -0.0783646, -0.11001797, -0.021044996, -0.06013344, -0.04063355, -0.09566213, -0.0027332064, -0.054325476, -0.012756522, -0.07795598, 0.009292462, -0.045779083, 0.0063116965, -0.059661258, 0.016208459, -0.036227033, 0.018023467, -0.042607244, 0.019224146, -0.026873393, 0.023964591, -0.027861275, 0.019463016, -0.018475424, 0.025666365, -0.015905868, 0.017893847, -0.011435829, 0.024489455, -0.006804505, 0.015300098, -0.005893507, 0.021564277, -0.00034539422, 0.01227663, -0.001805298, 0.017773021, 0.0038416486, 0.009244275, 0.0009852903, 0.013760047, 0.006195964, 0.0064746286, 0.0026938282, 0.009959627, 0.0071625044, 0.004119208, 0.00355482, 0.0066324025, 0.007150446, 0.0022388478, 0.0037941965, 0.003904212, 0.006509722, 0.0008306422, 0.0036123705, 0.0018030042, 0.005521167, -0.00014907392, 0.0031755941, 0.00029126342, 0.004396288, -0.00076632964, 0.0026134201, -0.00070733175},
		'{-0.040811576, -0.16744499, -0.0013990296, -0.24659619, -0.08905777, -0.12068868, -0.035101686, -0.18322004, -0.11222095, -0.0799173, -0.053682268, -0.12621841, -0.117192656, -0.046606373, -0.060886957, -0.0783646, -0.11001797, -0.021044996, -0.06013344, -0.04063355, -0.09566213, -0.0027332064, -0.054325476, -0.012756522, -0.07795598, 0.009292462, -0.045779083, 0.0063116965, -0.059661258, 0.016208459, -0.036227033, 0.018023467, -0.042607244, 0.019224146, -0.026873393, 0.023964591, -0.027861275, 0.019463016, -0.018475424, 0.025666365, -0.015905868, 0.017893847, -0.011435829, 0.024489455, -0.006804505, 0.015300098, -0.005893507, 0.021564277, -0.00034539422, 0.01227663, -0.001805298, 0.017773021, 0.0038416486, 0.009244275, 0.0009852903, 0.013760047, 0.006195964, 0.0064746286, 0.0026938282, 0.009959627, 0.0071625044, 0.004119208, 0.00355482, 0.0066324025, 0.007150446, 0.0022388478, 0.0037941965, 0.003904212, 0.006509722, 0.0008306422, 0.0036123705, 0.0018030042, 0.005521167, -0.00014907392, 0.0031755941, 0.00029126342, 0.004396288, -0.00076632964, 0.0026134201, -0.00070733175}};
	localparam real Ffi[0:3][0:79] = '{
		'{0.054977212, 0.27380404, -0.09682321, -0.13911411, 0.13286774, 0.14109056, -0.20146254, -0.06438994, 0.14257197, -0.013016365, -0.20590156, 0.016745165, 0.09660351, -0.12575768, -0.132206, 0.072398506, 0.025354939, -0.1647218, -0.026467597, 0.087769225, -0.03851404, -0.13279222, 0.064140536, 0.06664196, -0.07284027, -0.058710128, 0.10928026, 0.025568865, -0.07176878, 0.019808589, 0.10281957, -0.015350301, -0.044082917, 0.07231825, 0.059396178, -0.040833075, -0.0064497543, 0.085319765, 0.0040193177, -0.04499481, 0.024686437, 0.063301325, -0.039748963, -0.03132632, 0.03920768, 0.022798726, -0.058272038, -0.009166896, 0.035612084, -0.016647983, -0.05059351, 0.011176969, 0.019535823, -0.040521163, -0.025792554, 0.022519063, -4.7199166e-05, -0.04357123, 0.0027914792, 0.022744868, -0.014975273, -0.029587263, 0.02356174, 0.014402199, -0.020762067, -0.007838117, 0.030592768, 0.002643325, -0.01740584, 0.011695169, 0.024505815, -0.007320619, -0.008328141, 0.022224631, 0.010686009, -0.012184469, 0.0017177599, 0.021940462, -0.0038617796, -0.011335051},
		'{-0.054977212, -0.27380404, 0.09682321, 0.13911411, -0.13286774, -0.14109056, 0.20146254, 0.06438994, -0.14257197, 0.013016365, 0.20590156, -0.016745165, -0.09660351, 0.12575768, 0.132206, -0.072398506, -0.025354939, 0.1647218, 0.026467597, -0.087769225, 0.03851404, 0.13279222, -0.064140536, -0.06664196, 0.07284027, 0.058710128, -0.10928026, -0.025568865, 0.07176878, -0.019808589, -0.10281957, 0.015350301, 0.044082917, -0.07231825, -0.059396178, 0.040833075, 0.0064497543, -0.085319765, -0.0040193177, 0.04499481, -0.024686437, -0.063301325, 0.039748963, 0.03132632, -0.03920768, -0.022798726, 0.058272038, 0.009166896, -0.035612084, 0.016647983, 0.05059351, -0.011176969, -0.019535823, 0.040521163, 0.025792554, -0.022519063, 4.7199166e-05, 0.04357123, -0.0027914792, -0.022744868, 0.014975273, 0.029587263, -0.02356174, -0.014402199, 0.020762067, 0.007838117, -0.030592768, -0.002643325, 0.01740584, -0.011695169, -0.024505815, 0.007320619, 0.008328141, -0.022224631, -0.010686009, 0.012184469, -0.0017177599, -0.021940462, 0.0038617796, 0.011335051},
		'{0.2902459, -0.048090395, 0.1722119, -0.043068126, 0.21760303, -0.070462316, 0.13361703, -0.08219087, 0.1515946, -0.078621365, 0.096953146, -0.10009093, 0.09569856, -0.07691211, 0.06477738, -0.10274956, 0.051257875, -0.06900387, 0.03833797, -0.09536491, 0.01812269, -0.057806592, 0.017930374, -0.08217107, -0.004804195, -0.045484, 0.0032107749, -0.066406906, -0.01913248, -0.033528063, -0.0065455763, -0.050384194, -0.026659176, -0.02286643, -0.012244414, -0.035613447, -0.029142743, -0.01398146, -0.014827754, -0.022955867, -0.028161187, -0.0070262887, -0.0151775805, -0.012778579, -0.025036698, -0.0019286294, -0.014059162, -0.0050982754, -0.020809801, 0.0015224623, -0.012094923, 0.00029534003, -0.016247671, 0.0036084861, -0.009760273, 0.003740013, -0.01187366, 0.0046314257, -0.0073939264, 0.005625607, -0.008007896, 0.004879714, -0.0052166535, 0.0063410113, -0.004811392, 0.0046075317, -0.0033537855, 0.006240065, -0.0023285178, 0.004024518, -0.0018581408, 0.0056227297, -0.00052465417, 0.0032930924, -0.0007312022, 0.004727742, 0.0006825835, 0.0025309087, 5.8714853e-05, 0.003733309},
		'{-0.2902459, 0.048090395, -0.1722119, 0.043068126, -0.21760303, 0.070462316, -0.13361703, 0.08219087, -0.1515946, 0.078621365, -0.096953146, 0.10009093, -0.09569856, 0.07691211, -0.06477738, 0.10274956, -0.051257875, 0.06900387, -0.03833797, 0.09536491, -0.01812269, 0.057806592, -0.017930374, 0.08217107, 0.004804195, 0.045484, -0.0032107749, 0.066406906, 0.01913248, 0.033528063, 0.0065455763, 0.050384194, 0.026659176, 0.02286643, 0.012244414, 0.035613447, 0.029142743, 0.01398146, 0.014827754, 0.022955867, 0.028161187, 0.0070262887, 0.0151775805, 0.012778579, 0.025036698, 0.0019286294, 0.014059162, 0.0050982754, 0.020809801, -0.0015224623, 0.012094923, -0.00029534003, 0.016247671, -0.0036084861, 0.009760273, -0.003740013, 0.01187366, -0.0046314257, 0.0073939264, -0.005625607, 0.008007896, -0.004879714, 0.0052166535, -0.0063410113, 0.004811392, -0.0046075317, 0.0033537855, -0.006240065, 0.0023285178, -0.004024518, 0.0018581408, -0.0056227297, 0.00052465417, -0.0032930924, 0.0007312022, -0.004727742, -0.0006825835, -0.0025309087, -5.8714853e-05, -0.003733309}};
	localparam real Fbr[0:3][0:79] = '{
		'{-0.17863393, -0.09251931, 0.25321913, 0.060769558, -0.094903484, -0.20938554, 0.12451469, 0.11594125, 0.0045285556, -0.22019, -0.020327035, 0.11464327, 0.07871964, -0.14600335, -0.12326026, 0.07073361, 0.10587191, -0.03472484, -0.15567382, 0.01074123, 0.08695919, 0.06320277, -0.12213215, -0.03906609, 0.039970078, 0.114279784, -0.050810527, -0.062453806, -0.010855579, 0.11047875, 0.022644024, -0.056922436, -0.045581665, 0.06621784, 0.07022722, -0.031390827, -0.05502016, 0.0076479567, 0.08025168, -0.00015333144, -0.041625693, -0.03991569, 0.05785849, 0.0237445, -0.015819622, -0.06127297, 0.019107524, 0.033094063, 0.009797943, -0.054634042, -0.017620465, 0.027840206, 0.025681186, -0.029113853, -0.039054655, 0.0134079205, 0.028188987, 0.0012624935, -0.0407923, -0.002626315, 0.019549819, 0.023973053, -0.026847044, -0.013880414, 0.00563754, 0.03233093, -0.0061533004, -0.017273117, -0.0070908256, 0.026605913, 0.011943759, -0.013395881, -0.014150508, 0.0122761205, 0.021284029, -0.005421758, -0.01424092, -0.0032561799, 0.020444404, 0.0026938305},
		'{-0.17863393, -0.09251931, 0.25321913, 0.060769558, -0.094903484, -0.20938554, 0.12451469, 0.11594125, 0.0045285556, -0.22019, -0.020327035, 0.11464327, 0.07871964, -0.14600335, -0.12326026, 0.07073361, 0.10587191, -0.03472484, -0.15567382, 0.01074123, 0.08695919, 0.06320277, -0.12213215, -0.03906609, 0.039970078, 0.114279784, -0.050810527, -0.062453806, -0.010855579, 0.11047875, 0.022644024, -0.056922436, -0.045581665, 0.06621784, 0.07022722, -0.031390827, -0.05502016, 0.0076479567, 0.08025168, -0.00015333144, -0.041625693, -0.03991569, 0.05785849, 0.0237445, -0.015819622, -0.06127297, 0.019107524, 0.033094063, 0.009797943, -0.054634042, -0.017620465, 0.027840206, 0.025681186, -0.029113853, -0.039054655, 0.0134079205, 0.028188987, 0.0012624935, -0.0407923, -0.002626315, 0.019549819, 0.023973053, -0.026847044, -0.013880414, 0.00563754, 0.03233093, -0.0061533004, -0.017273117, -0.0070908256, 0.026605913, 0.011943759, -0.013395881, -0.014150508, 0.0122761205, 0.021284029, -0.005421758, -0.01424092, -0.0032561799, 0.020444404, 0.0026938305},
		'{-0.040811576, 0.16744499, -0.0013990296, 0.24659619, -0.08905777, 0.12068868, -0.035101686, 0.18322004, -0.11222095, 0.0799173, -0.053682268, 0.12621841, -0.117192656, 0.046606373, -0.060886957, 0.0783646, -0.11001797, 0.021044996, -0.06013344, 0.04063355, -0.09566213, 0.0027332064, -0.054325476, 0.012756522, -0.07795598, -0.009292462, -0.045779083, -0.0063116965, -0.059661258, -0.016208459, -0.036227033, -0.018023467, -0.042607244, -0.019224146, -0.026873393, -0.023964591, -0.027861275, -0.019463016, -0.018475424, -0.025666365, -0.015905868, -0.017893847, -0.011435829, -0.024489455, -0.006804505, -0.015300098, -0.005893507, -0.021564277, -0.00034539422, -0.01227663, -0.001805298, -0.017773021, 0.0038416486, -0.009244275, 0.0009852903, -0.013760047, 0.006195964, -0.0064746286, 0.0026938282, -0.009959627, 0.0071625044, -0.004119208, 0.00355482, -0.0066324025, 0.007150446, -0.0022388478, 0.0037941965, -0.003904212, 0.006509722, -0.0008306422, 0.0036123705, -0.0018030042, 0.005521167, 0.00014907392, 0.0031755941, -0.00029126342, 0.004396288, 0.00076632964, 0.0026134201, 0.00070733175},
		'{-0.040811576, 0.16744499, -0.0013990296, 0.24659619, -0.08905777, 0.12068868, -0.035101686, 0.18322004, -0.11222095, 0.0799173, -0.053682268, 0.12621841, -0.117192656, 0.046606373, -0.060886957, 0.0783646, -0.11001797, 0.021044996, -0.06013344, 0.04063355, -0.09566213, 0.0027332064, -0.054325476, 0.012756522, -0.07795598, -0.009292462, -0.045779083, -0.0063116965, -0.059661258, -0.016208459, -0.036227033, -0.018023467, -0.042607244, -0.019224146, -0.026873393, -0.023964591, -0.027861275, -0.019463016, -0.018475424, -0.025666365, -0.015905868, -0.017893847, -0.011435829, -0.024489455, -0.006804505, -0.015300098, -0.005893507, -0.021564277, -0.00034539422, -0.01227663, -0.001805298, -0.017773021, 0.0038416486, -0.009244275, 0.0009852903, -0.013760047, 0.006195964, -0.0064746286, 0.0026938282, -0.009959627, 0.0071625044, -0.004119208, 0.00355482, -0.0066324025, 0.007150446, -0.0022388478, 0.0037941965, -0.003904212, 0.006509722, -0.0008306422, 0.0036123705, -0.0018030042, 0.005521167, 0.00014907392, 0.0031755941, -0.00029126342, 0.004396288, 0.00076632964, 0.0026134201, 0.00070733175}};
	localparam real Fbi[0:3][0:79] = '{
		'{-0.054977212, 0.27380404, 0.09682321, -0.13911411, -0.13286774, 0.14109056, 0.20146254, -0.06438994, -0.14257197, -0.013016365, 0.20590156, 0.016745165, -0.09660351, -0.12575768, 0.132206, 0.072398506, -0.025354939, -0.1647218, 0.026467597, 0.087769225, 0.03851404, -0.13279222, -0.064140536, 0.06664196, 0.07284027, -0.058710128, -0.10928026, 0.025568865, 0.07176878, 0.019808589, -0.10281957, -0.015350301, 0.044082917, 0.07231825, -0.059396178, -0.040833075, 0.0064497543, 0.085319765, -0.0040193177, -0.04499481, -0.024686437, 0.063301325, 0.039748963, -0.03132632, -0.03920768, 0.022798726, 0.058272038, -0.009166896, -0.035612084, -0.016647983, 0.05059351, 0.011176969, -0.019535823, -0.040521163, 0.025792554, 0.022519063, 4.7199166e-05, -0.04357123, -0.0027914792, 0.022744868, 0.014975273, -0.029587263, -0.02356174, 0.014402199, 0.020762067, -0.007838117, -0.030592768, 0.002643325, 0.01740584, 0.011695169, -0.024505815, -0.007320619, 0.008328141, 0.022224631, -0.010686009, -0.012184469, -0.0017177599, 0.021940462, 0.0038617796, -0.011335051},
		'{0.054977212, -0.27380404, -0.09682321, 0.13911411, 0.13286774, -0.14109056, -0.20146254, 0.06438994, 0.14257197, 0.013016365, -0.20590156, -0.016745165, 0.09660351, 0.12575768, -0.132206, -0.072398506, 0.025354939, 0.1647218, -0.026467597, -0.087769225, -0.03851404, 0.13279222, 0.064140536, -0.06664196, -0.07284027, 0.058710128, 0.10928026, -0.025568865, -0.07176878, -0.019808589, 0.10281957, 0.015350301, -0.044082917, -0.07231825, 0.059396178, 0.040833075, -0.0064497543, -0.085319765, 0.0040193177, 0.04499481, 0.024686437, -0.063301325, -0.039748963, 0.03132632, 0.03920768, -0.022798726, -0.058272038, 0.009166896, 0.035612084, 0.016647983, -0.05059351, -0.011176969, 0.019535823, 0.040521163, -0.025792554, -0.022519063, -4.7199166e-05, 0.04357123, 0.0027914792, -0.022744868, -0.014975273, 0.029587263, 0.02356174, -0.014402199, -0.020762067, 0.007838117, 0.030592768, -0.002643325, -0.01740584, -0.011695169, 0.024505815, 0.007320619, -0.008328141, -0.022224631, 0.010686009, 0.012184469, 0.0017177599, -0.021940462, -0.0038617796, 0.011335051},
		'{0.2902459, 0.048090395, 0.1722119, 0.043068126, 0.21760303, 0.070462316, 0.13361703, 0.08219087, 0.1515946, 0.078621365, 0.096953146, 0.10009093, 0.09569856, 0.07691211, 0.06477738, 0.10274956, 0.051257875, 0.06900387, 0.03833797, 0.09536491, 0.01812269, 0.057806592, 0.017930374, 0.08217107, -0.004804195, 0.045484, 0.0032107749, 0.066406906, -0.01913248, 0.033528063, -0.0065455763, 0.050384194, -0.026659176, 0.02286643, -0.012244414, 0.035613447, -0.029142743, 0.01398146, -0.014827754, 0.022955867, -0.028161187, 0.0070262887, -0.0151775805, 0.012778579, -0.025036698, 0.0019286294, -0.014059162, 0.0050982754, -0.020809801, -0.0015224623, -0.012094923, -0.00029534003, -0.016247671, -0.0036084861, -0.009760273, -0.003740013, -0.01187366, -0.0046314257, -0.0073939264, -0.005625607, -0.008007896, -0.004879714, -0.0052166535, -0.0063410113, -0.004811392, -0.0046075317, -0.0033537855, -0.006240065, -0.0023285178, -0.004024518, -0.0018581408, -0.0056227297, -0.00052465417, -0.0032930924, -0.0007312022, -0.004727742, 0.0006825835, -0.0025309087, 5.8714853e-05, -0.003733309},
		'{-0.2902459, -0.048090395, -0.1722119, -0.043068126, -0.21760303, -0.070462316, -0.13361703, -0.08219087, -0.1515946, -0.078621365, -0.096953146, -0.10009093, -0.09569856, -0.07691211, -0.06477738, -0.10274956, -0.051257875, -0.06900387, -0.03833797, -0.09536491, -0.01812269, -0.057806592, -0.017930374, -0.08217107, 0.004804195, -0.045484, -0.0032107749, -0.066406906, 0.01913248, -0.033528063, 0.0065455763, -0.050384194, 0.026659176, -0.02286643, 0.012244414, -0.035613447, 0.029142743, -0.01398146, 0.014827754, -0.022955867, 0.028161187, -0.0070262887, 0.0151775805, -0.012778579, 0.025036698, -0.0019286294, 0.014059162, -0.0050982754, 0.020809801, 0.0015224623, 0.012094923, 0.00029534003, 0.016247671, 0.0036084861, 0.009760273, 0.003740013, 0.01187366, 0.0046314257, 0.0073939264, 0.005625607, 0.008007896, 0.004879714, 0.0052166535, 0.0063410113, 0.004811392, 0.0046075317, 0.0033537855, 0.006240065, 0.0023285178, 0.004024518, 0.0018581408, 0.0056227297, 0.00052465417, 0.0032930924, 0.0007312022, 0.004727742, -0.0006825835, 0.0025309087, -5.8714853e-05, 0.003733309}};
	localparam real hf[0:1199] = {0.23903719, -0.056577254, -0.046376806, 0.009240281, 0.16428359, -0.13344508, -0.0036647443, 0.01928589, 0.081619464, -0.15000962, 0.05185026, 0.011636511, 0.014241237, -0.11663765, 0.09115172, -0.010857091, -0.024764504, -0.05822209, 0.098571725, -0.037874848, -0.034566384, -0.0019830666, 0.07477467, -0.058038898, -0.023895573, 0.032810993, 0.03275979, -0.064085096, -0.0055858963, 0.03981509, -0.009921085, -0.055135515, 0.009022917, 0.024662416, -0.03888094, -0.035908896, 0.013744869, -0.00015487392, -0.04764395, -0.013902288, 0.008398102, -0.021689452, -0.03832304, 0.0039017962, -0.0027806722, -0.031541757, -0.018921323, 0.0134365605, -0.013971439, -0.027936192, 0.00094403164, 0.014351925, -0.020490887, -0.01479963, 0.013927031, 0.009275766, -0.020404473, 0.0010919541, 0.017087722, 0.0021609426, -0.014691741, 0.013364744, 0.01189166, -0.003458948, -0.006250252, 0.018378805, 0.0025779814, -0.0056395885, 0.0016081632, 0.015981153, -0.0061094626, -0.004325947, 0.0064796824, 0.008769799, -0.010830792, -0.00087981566, 0.007551678, 0.0004959182, -0.010572402, 0.0028033704, 0.0055375565, -0.0055937036, -0.0064739278, 0.0051599727, 0.0020609503, -0.0078387195, -0.00088632095, 0.005486435, -0.0011527935, -0.0064021344, 0.0038024418, 0.0040134266, -0.0029316158, -0.002772526, 0.0060780346, 0.0016068702, -0.0029507598, 0.0011090921, 0.0056674257, -0.0007025566, -0.001641975, 0.0036829025, 0.003353879, -0.0021434487, 0.00015665147, 0.004262454, 0.00043916042, -0.0024323983, 0.0016177294, 0.0030825865, -0.001862258, -0.0017671462, 0.0022367118, 0.0009908297, -0.0028540406, -0.00064182235, 0.0019474562, -0.0010174464, -0.0024938714, 0.00040492573, 0.0010448572, -0.0022089037, -0.0012531686, 0.0009990553, -1.0437184e-05, -0.0023265942, 0.00018164712, 0.001029527, -0.0008038651, -0.0015748176, 0.0012171555, 0.0006254468, -0.0011118401, -0.00043450092, 0.0015528711, 4.9232138e-05, -0.00094108394, 0.00058160716, 0.0012239799, -0.0004343547, -0.0004725073, 0.001127973, 0.0005082042, -0.0006586299, 4.6858797e-05, 0.0011158069, -0.0002360883, -0.0005945838, 0.00041119408, 0.00068544026, -0.0007235973, -0.00032931016, 0.0005225105, 9.9579425e-05, -0.0008319858, -5.902313e-06, 0.00040127503, -0.0003839079, -0.00060940516, 0.00024349481, 0.00015031172, -0.00060723675, -0.00021633696, 0.00034474264, -0.00010345545, -0.00054791843, 0.00016091713, 0.00029593165, -0.0002623835, -0.0002949932, 0.000385986, 0.000151193, -0.00028780816, 1.084417e-05, 0.00041159766, -1.26556315e-05, -0.00020057078, 0.00024225442, 0.00027615347, -0.00013008782, -5.9104073e-05, 0.00032984538, 6.906533e-05, -0.00016860482, 7.138953e-05, 0.00027448742, -0.00011477901, -0.00013299152, 0.0001450063, 0.0001303883, -0.00021180927, -5.463472e-05, 0.00014781408, -2.7808315e-05, -0.0002061253, 2.6564689e-05, 9.555136e-05, -0.00013779633, -0.0001241317, 7.916516e-05, 2.0756184e-05, -0.00017001014, -1.4608162e-05, 8.995813e-05, -4.3355023e-05, -0.00013094475, 7.487308e-05, 6.459199e-05, -7.5454125e-05, -5.2193198e-05, 0.000115488736, 2.0983176e-05, -7.1249924e-05, 2.7314725e-05, 0.00010352842, -2.030821e-05, -4.1046686e-05, 7.761436e-05, 5.584598e-05, -4.4414155e-05, -2.4226397e-06, 8.679232e-05, -1.3141753e-06, -4.638906e-05, 2.807657e-05, 6.116444e-05, -4.4363027e-05, -3.0722178e-05, 4.088765e-05, 1.8588575e-05, -6.0568334e-05, -7.4315167e-06, 3.535451e-05, -2.095851e-05, -5.0250837e-05, 1.29890805e-05, 1.7861572e-05, -4.3364787e-05, -2.3574563e-05, 2.3606332e-05, -2.2271104e-06, -4.4279313e-05, 5.587432e-06, 2.2796748e-05, -1.6782578e-05, -2.8430753e-05, 2.5723135e-05, 1.3595162e-05, -2.1664937e-05, -5.707431e-06, 3.143047e-05, 1.4546162e-06, -1.7331313e-05, 1.3766452e-05, 2.3991272e-05, -8.367861e-06, -7.57829e-06, 2.3477261e-05, 9.307361e-06, -1.2732551e-05, 2.668597e-06, 2.2106002e-05, -5.4039187e-06, -1.1290444e-05, 9.465061e-06, 1.2792604e-05, -1.46239e-05, -5.9522877e-06, 1.1091634e-05, 9.051408e-07, -1.6196838e-05, 3.626266e-07, 8.170177e-06, -8.496937e-06, -1.1340891e-05, 5.0589033e-06, 2.8765296e-06, -1.2483393e-05, -3.39326e-06, 6.7605965e-06, -2.2419993e-06, -1.08456625e-05, 3.9409356e-06, 5.538049e-06, -5.3080794e-06, -5.5301907e-06, 8.0629225e-06, 2.539449e-06, -5.6583185e-06, 6.0073427e-07, 8.191286e-06, -6.9399124e-07, -3.8039354e-06, 5.0575104e-06, 5.2242754e-06, -2.8979214e-06, -9.610125e-07, 6.567052e-06, 1.0058891e-06, -3.492535e-06, 1.5718692e-06, 5.261336e-06, -2.5883094e-06, -2.6374971e-06, 2.919471e-06, 2.2952581e-06, -4.3607315e-06, -9.970679e-07, 2.857432e-06, -8.2797925e-07, -4.0794885e-06, 6.280356e-07, 1.7422229e-06, -2.9021387e-06, -2.3364687e-06, 1.6326735e-06, 2.402107e-07, -3.399242e-06, -1.3064476e-07, 1.7874688e-06, -9.951585e-07, -2.5066513e-06, 1.6023358e-06, 1.2356509e-06, -1.5649143e-06, -8.875635e-07, 2.3254472e-06, 3.511592e-07, -1.4136614e-06, 6.799244e-07, 2.0069417e-06, -4.560163e-07, -7.6896475e-07, 1.621302e-06, 1.0125854e-06, -9.0188763e-07, 1.0838011e-08, 1.7325017e-06, -1.254113e-07, -9.0496854e-07, 6.017416e-07, 1.1685662e-06, -9.4705706e-07, -5.688418e-07, 8.2722744e-07, 3.0056216e-07, -1.219693e-06, -9.9564744e-08, 6.8940943e-07, -4.7449282e-07, -9.712672e-07, 2.957343e-07, 3.2593118e-07, -8.884072e-07, -4.1816645e-07, 4.8665123e-07, -7.3665895e-08, -8.7171094e-07, 1.6041015e-07, 4.5015815e-07, -3.5119737e-07, -5.326038e-07, 5.418449e-07, 2.5379984e-07, -4.3163485e-07, -7.437376e-08, 6.3004137e-07, 8.962163e-09, -3.3150576e-07, 3.0322713e-07, 4.6143782e-07, -1.8120618e-07, -1.310274e-07, 4.7792867e-07, 1.5998009e-07, -2.58456e-07, 7.100539e-08, 4.32371e-07, -1.3000246e-07, -2.2060979e-07, 1.986052e-07, 2.3576192e-07, -3.026566e-07, -1.0909697e-07, 2.2163921e-07, -2.5306413e-09, -3.2112217e-07, 1.6883664e-08, 1.5625234e-07, -1.8343192e-07, -2.1499358e-07, 1.0673519e-07, 4.786528e-08, -2.528132e-07, -5.3503456e-08, 1.3536831e-07, -5.2761305e-08, -2.1111244e-07, 8.978269e-08, 1.06554204e-07, -1.097939e-07, -1.0024878e-07, 1.6553369e-07, 4.4678764e-08, -1.1220572e-07, 2.189342e-08, 1.613825e-07, -1.9268386e-08, -7.203007e-08, 1.0691534e-07, 9.7803216e-08, -6.085932e-08, -1.439441e-08, 1.3177639e-07, 1.2669572e-08, -6.981926e-08, 3.498757e-08, 1.01415e-07, -5.704394e-08, -5.052182e-08, 5.9581375e-08, 4.027415e-08, -8.889118e-08, -1.6883131e-08, 5.604816e-08, -2.1468104e-08, -7.991713e-08, 1.5107494e-08, 3.2369986e-08, -6.055461e-08, -4.3148642e-08, 3.3864257e-08, 2.18074e-09, -6.771711e-08, 1.0669722e-09, 3.549939e-08, -2.1676367e-08, -4.7833446e-08, 3.441283e-08, 2.345563e-08, -3.1769744e-08, -1.4751694e-08, 4.697896e-08, 5.4814357e-09, -2.7580162e-08, 1.601829e-08, 3.89815e-08, -1.0289445e-08, -1.4058324e-08, 3.3504808e-08, 1.828389e-08, -1.8474266e-08, 1.5237563e-09, 3.4307146e-08, -4.3578865e-09, -1.7804986e-08, 1.2844849e-08, 2.2075891e-08, -2.0006997e-08, -1.0628623e-08, 1.6675804e-08, 4.4765187e-09, -2.4460686e-08, -1.1725421e-09, 1.3356231e-08, -1.0631065e-08, -1.8702641e-08, 6.483426e-09, 5.8222533e-09, -1.8181064e-08, -7.306587e-09, 9.8994235e-09, -2.1075506e-09, -1.7136626e-08, 4.126109e-09, 8.800645e-09, -7.3706787e-09, -9.923937e-09, 1.1306756e-08, 4.6675335e-09, -8.628178e-09, -7.0388245e-10, 1.2554064e-08, -2.3408422e-10, -6.3577685e-09, 6.596456e-09, 8.806126e-09, -3.8872323e-09, -2.2448061e-09, 9.698616e-09, 2.6489575e-09, -5.219948e-09, 1.7346367e-09, 8.435354e-09, -3.0418588e-09, -4.28281e-09, 4.122399e-09, 4.313317e-09, -6.2462773e-09, -1.9641828e-09, 4.401484e-09, -4.473801e-10, -6.3534378e-09, 5.407512e-10, 2.9667435e-09, -3.913248e-09, -4.056658e-09, 2.2500861e-09, 7.611298e-10, -5.093392e-09, -7.850426e-10, 2.7122853e-09, -1.2071054e-09, -4.0872674e-09, 2.0057669e-09, 2.0496311e-09, -2.2573325e-09, -1.7892504e-09, 3.3848249e-09, 7.765635e-10, -2.2137703e-09, 6.344276e-10, 3.170153e-09, -4.85774e-10, -1.3517434e-09, 2.246657e-09, 1.8195114e-09, -1.2673408e-09, -1.8778726e-10, 2.6360196e-09, 1.0753591e-10, -1.3893875e-09, 7.708468e-10, 1.9463269e-09, -1.2392986e-09, -9.623969e-10, 1.2138925e-09, 6.9130207e-10, -1.8032444e-09, -2.7623248e-10, 1.097577e-09, -5.253384e-10, -1.558567e-09, 3.5085534e-10, 5.979019e-10, -1.2572086e-09, -7.883495e-10, 6.980945e-10, -7.28967e-12, -1.3451111e-09, 9.4612825e-11, 7.0175876e-10, -4.664454e-10, -9.086293e-10, 7.3306694e-10, 4.4183632e-10, -6.4225203e-10, -2.3534305e-10, 9.458945e-10, 7.80528e-11, -5.3598964e-10, 3.6661402e-10, 7.5420803e-10, -2.2880702e-10, -2.5423344e-10, 6.8877803e-10, 3.2555897e-10, -3.7734316e-10, 5.5978822e-11, 6.767958e-10, -1.2346603e-10, -3.4943906e-10, 2.7177485e-10, 4.1427922e-10, -4.1994003e-10, -1.9732237e-10, 3.3472522e-10, 5.883345e-11, -4.8899595e-10, -7.354714e-12, 2.5745744e-10, -2.3446747e-10, -3.58634e-10, 1.4038243e-10, 1.0210227e-10, -3.7053643e-10, -1.2488001e-10, 2.0058077e-10, -5.4688632e-11, -3.3566602e-10, 1.002722e-10, 1.71433e-10, -1.5387734e-10, -1.8338935e-10, 2.3456928e-10, 8.500832e-11, -1.7197076e-10, 1.4837351e-12, 2.49249e-10, -1.2775306e-11, -1.213987e-10, 1.420233e-10, 1.6714122e-10, -8.262086e-11, -3.735388e-11, 1.9611368e-10, 4.190402e-11, -1.0499606e-10, 4.0773388e-11, 1.6397626e-10, -6.9364424e-11, -8.2765364e-11, 8.513583e-11, 7.8061155e-11, -1.2831633e-10, -3.481403e-11, 8.712096e-11, -1.6732995e-11, -1.2527049e-10, 1.4815689e-11, 5.6020587e-11, -8.281549e-11, -7.60483e-11, 4.7146446e-11, 1.1312403e-11, -1.0224596e-10, -1.00117145e-11, 5.4170977e-11, -2.7043843e-11, -7.8797455e-11, 4.4135452e-11, 3.9252043e-11, -4.6192872e-11, -3.1402166e-11, 6.893752e-11, 1.3171089e-11, -4.351415e-11, 1.652589e-11, 6.205828e-11, -1.1664765e-11, -2.5179353e-11, 4.691772e-11, 3.3575264e-11, -2.6252545e-11, -1.7598609e-12, 5.2548122e-11, -7.3253437e-13, -2.7557769e-11, 1.6772701e-11, 3.7172775e-11, -2.6641982e-11, -1.8237111e-11, 2.4637521e-11, 1.1521935e-11, -3.6442085e-11, -4.296168e-12, 2.1416377e-11, -1.2368233e-11, -3.0278686e-11, 7.951902e-12, 1.0940336e-11, -2.5970887e-11, -1.4239348e-11, 1.4322662e-11, -1.1507129e-12, -2.662969e-11, 3.332645e-12, 1.38228404e-11, -9.947803e-12, -1.7163118e-11, 1.5495927e-11, 8.2665185e-12, -1.2937575e-11, -3.512875e-12, 1.8977715e-11, 9.312016e-13, -1.0375924e-11, 8.220096e-12, 1.4530316e-11, -5.0157166e-12, -4.536437e-12, 1.4097329e-11, 5.6963457e-12, -7.676661e-12, 1.6185608e-12, 1.33052085e-11, -3.1782758e-12, -6.8335754e-12, 5.7101086e-12, 7.719588e-12, -8.761526e-12, -3.631843e-12, 6.695079e-12, 5.666634e-13, -9.742602e-12, 1.7137145e-13, 4.9403693e-12, -5.104583e-12, -6.8440167e-12, 3.0098257e-12, 1.7516496e-12, -7.5218685e-12, -2.0696214e-12, 4.0493425e-12, -1.3377434e-12, -6.5507734e-12, 2.3489977e-12, 3.326747e-12, -3.194753e-12, -3.3572195e-12, 4.841889e-12, 1.5298277e-12, -3.416e-12, 3.3694139e-13, 4.931802e-12, -4.1430165e-13, -2.3060056e-12, 3.0301805e-12, 3.1541033e-12, -1.7429572e-12, -5.9555876e-13, 3.951248e-12, 6.1656274e-13, -2.1044746e-12, 9.328125e-13, 3.174976e-12, -1.5509085e-12, -1.5925316e-12, 1.7500467e-12, 1.3939086e-12, -2.6245063e-12, -6.056207e-13, 1.7185936e-12, -4.8723834e-13, -2.4613378e-12, 3.7431505e-13, 1.0511981e-12, -1.7405205e-12, -1.4153557e-12, 9.820685e-13, 1.4830509e-13, -2.045425e-12, -8.719608e-14, 1.078248e-12, -5.963031e-13, -1.5123815e-12, 9.590977e-13, 7.479879e-13, -9.413492e-13, -5.3937237e-13, 1.3985704e-12, 2.1590919e-13, -8.522749e-13, 4.0515228e-13, 1.2103922e-12, -2.710028e-13, -4.652271e-13, 9.743356e-13, 6.1363984e-13, -5.4115816e-13, 4.3346716e-15, 1.0439734e-12, -7.152961e-14, -5.447469e-13, 3.6108096e-13, 7.0628827e-13, -5.676717e-13, -3.4354876e-13, 4.9817133e-13, 1.8415388e-13, -7.338075e-13, -6.138003e-14, 4.1629802e-13, -2.8328034e-13, -5.858864e-13, 1.7694975e-13, 1.9796273e-13, -5.339739e-13, -2.5365465e-13, 2.9259809e-13, -4.2781947e-14, -5.25399e-13, 9.4865074e-14, 2.7132075e-13, -2.1050177e-13, -3.2216084e-13, 3.2534034e-13, 1.5350748e-13, -2.5969976e-13, -4.644219e-14, 3.7944105e-13, 6.1238496e-15, -2.0002373e-13, 1.8137262e-13, 2.786792e-13, -1.08651776e-13, -7.959608e-14, 2.8734014e-13, 9.744862e-14, -1.5557243e-13, 4.21126e-14, 2.6064283e-13, -7.7348264e-14, -1.3314051e-13, 1.1923485e-13, 1.426905e-13, -1.8179619e-13, -6.617664e-14, 1.3345648e-13, -7.496745e-16, -1.9345163e-13, 9.704703e-15, 9.4348276e-14, -1.0994244e-13, -1.2992451e-13, 6.398412e-14, 2.9179733e-14, -1.5211905e-13, -3.280078e-14, 8.145635e-14, -3.1480864e-14, -1.2735936e-13, 5.36036e-14, 6.429631e-14, -6.599147e-14, -6.0783206e-14, 9.9479744e-14, 2.7129146e-14, -6.7624685e-14, 1.2783077e-14, 9.725011e-14, -1.1393148e-14, -4.355447e-14, 6.414319e-14, 5.91409e-14, -3.652807e-14, -8.878608e-15, 7.9327875e-14, 7.915383e-15, -4.2035992e-14, 2.0909867e-14, 6.1218805e-14, -3.4143166e-14, -3.0502605e-14, 3.5816368e-14, 2.4479474e-14, -5.346002e-14, -1.0281065e-14, 3.378441e-14, -1.2724337e-14, -4.8188782e-14, 9.000922e-15, 1.958574e-14, -3.6354637e-14, -2.6125325e-14, 2.0347237e-14, 1.4170076e-15, -4.077916e-14, 4.9403117e-16, 2.1389334e-14, -1.2979838e-14, -2.8889444e-14, 2.0624947e-14, 1.4177127e-14, -1.910823e-14, -8.999874e-15, 2.8267477e-14, 3.365282e-15, -1.663186e-14, 9.549115e-15, 2.3517741e-14, -6.1461697e-15, -8.5154204e-15, 2.013078e-14, 1.1088403e-14, -1.1104357e-14, 8.6695934e-16, 2.067033e-14, -2.5488255e-15, -1.07312984e-14, 7.703018e-15, 1.33437556e-14, -1.2002541e-14, -6.429101e-15, 1.0036511e-14, 2.756614e-15, -1.4724213e-14, -7.3880294e-16, 8.060058e-15, -6.3554767e-15, -1.1289081e-14, 3.8806133e-15, 3.5341842e-15, -1.0930514e-14, -4.4410945e-15, 5.953361e-15, -1.2430522e-15, -1.0330117e-14, 2.4478962e-15, 5.306518e-15, -4.4236728e-15, -6.004606e-15, 6.789148e-15, 2.8262453e-15, -5.195027e-15, -4.5543326e-16, 7.560731e-15, -1.2475899e-16, -3.8388605e-15, 3.950191e-15, 5.3190895e-15, -2.3302567e-15, -1.3666794e-15, 5.8337247e-15, 1.6169612e-15, -3.1411114e-15, 1.031731e-15, 5.0872625e-15, -1.8138419e-15, -2.5840159e-15, 2.4759461e-15, 2.613043e-15, -3.7531793e-15, -1.1914624e-15, 2.651249e-15, -2.535249e-16, -3.8282006e-15, 3.1738145e-16, 1.792491e-15, -2.3463746e-15, -2.4522919e-15, 1.3501114e-15, 4.6603213e-16, -3.0652225e-15, -4.841344e-16, 1.6328483e-15, -7.2078856e-16, -2.4663181e-15, 1.1992071e-15, 1.2373428e-15, -1.3567271e-15, -1.0859185e-15, 2.0349842e-15, 4.7226894e-16, -1.3341564e-15, 3.7413691e-16, 1.9110107e-15, -2.884382e-16, -8.174619e-16, 1.348384e-15, 1.1009686e-15, -7.610265e-16, -1.1708761e-16, 1.5871335e-15, 7.057515e-17, -8.367997e-16, 4.612715e-16, 1.1751712e-15, -7.4224137e-16, -5.813567e-16, 7.299883e-16, 4.2081267e-16, -1.084709e-15, -1.6876016e-16, 6.617867e-16, -3.1245285e-16, -9.399971e-16, 2.0931193e-16, 3.61982e-16, -7.551073e-16, -4.7764606e-16, 4.19496e-16, -2.343996e-18, -8.10251e-16, 5.403633e-17, 4.2286145e-16, -2.7951973e-16, -5.4900266e-16, 4.3958625e-16, 2.6712314e-16, -3.8641609e-16, -1.4408786e-16, 5.692695e-16, 4.8260844e-17, -3.2333656e-16, 2.1888496e-16, 4.5512605e-16, -1.3684209e-16, -1.5414671e-16, 4.1396144e-16, 1.9762617e-16, -2.2688286e-16, 3.2686786e-17, 4.0786873e-16, -7.288289e-17, -2.1066367e-16, 1.6304098e-16, 2.5052482e-16, -2.5204995e-16, -1.1941897e-16, 2.0148946e-16, 3.665104e-17, -2.9443006e-16, -5.0741794e-18, 1.5540163e-16, -1.402983e-16, -2.1654863e-16, 8.409328e-17, 6.2049676e-17, -2.2282234e-16, -7.604021e-17, 1.2066377e-16, -3.2426003e-17, -2.0238655e-16, 5.966288e-17, 1.034014e-16, -9.239042e-17, -1.1102243e-16, 1.4089534e-16, 5.1516355e-17, -1.03566977e-16, 2.7007362e-19, 1.5014484e-16, -7.3684595e-18, -7.3324506e-17, 8.51073e-17, 1.0099427e-16, -4.9550762e-17, -2.279296e-17, 1.1799334e-16, 2.5673345e-17, -6.319392e-17, 2.4305675e-17, 9.891874e-17, -4.1422856e-17, -4.9948434e-17, 5.1151986e-17, 4.7328767e-17, -7.7123124e-17, -2.114028e-17, 5.249128e-17, -9.763135e-18, -7.549693e-17, 8.76037e-18, 3.3862246e-17, -4.9680593e-17, -4.5992003e-17, 2.8300896e-17, 6.9675665e-18, -6.154662e-17, -6.2558297e-18, 3.261919e-17, -1.616688e-17, -4.756153e-17, 2.6412777e-17, 2.3703251e-17, -2.7770667e-17, -1.9082496e-17, 4.1457267e-17, 8.02482e-18, -2.6230152e-17, 9.796596e-18, 3.7418835e-17, -6.945198e-18, -1.5234642e-17, 2.8169536e-17, 2.0328207e-17, -1.5770227e-17, -1.1394802e-18, 3.164591e-17, -3.2562355e-19, -1.6601574e-17, 1.0044521e-17, 2.2451783e-17, -1.5966703e-17, -1.1020921e-17, 1.481977e-17, 7.029552e-18, -2.19265e-17, -2.6358658e-18, 1.2916152e-17, -7.372336e-18, -1.826638e-17, 4.7503903e-18, 6.6278893e-18, -1.5603859e-17, -8.634589e-18, 8.609169e-18, -6.525927e-19, -1.6044528e-17, 1.9489192e-18, 8.331167e-18, -5.964738e-18, -1.037425e-17, 9.296625e-18, 5.000055e-18, -7.785942e-18, -2.1628883e-18, 1.1424007e-17, 5.858807e-19, -6.2610566e-18, 4.913737e-18, 8.770813e-18, -3.0023494e-18, -2.753312e-18, 8.4750535e-18, 3.4623657e-18, -4.6168925e-18, 9.545539e-19, 8.020238e-18, -1.8852435e-18, -4.120683e-18, 3.427037e-18, 4.670584e-18, -5.2607545e-18, -2.1993144e-18, 4.0310525e-18, 3.6560315e-19, -5.867471e-18, 9.043013e-20, 2.9829303e-18, -3.056825e-18, -4.133909e-18, 1.8041068e-18, 1.0662837e-18, -4.5244348e-18, -1.2632435e-18, 2.436579e-18, -7.9568426e-19, -3.9506986e-18, 1.4005668e-18, 2.0070983e-18, -1.918856e-18, -2.0337993e-18, 2.9092536e-18, 9.27921e-19, -2.0576966e-18, 1.9057048e-19, 2.9715436e-18, -2.4309225e-19, -1.3933192e-18, 1.8168635e-18, 1.9066255e-18, -1.045802e-18, -3.6464952e-19, 2.377869e-18, 3.8009696e-19, -1.266912e-18, 5.5694417e-19, 1.9158241e-18, -9.272453e-19, -9.613686e-19, 1.0518002e-18, 8.459643e-19, -1.5778744e-18, -3.682704e-19, 1.0357111e-18, -2.8725574e-19, -1.4837246e-18, 2.2225118e-19, 6.3569233e-19, -1.0445882e-18, -8.5640713e-19, 5.897324e-19, 9.2414066e-20, -1.2315208e-18, -5.70255e-20, 6.4941547e-19, -3.568125e-19, -9.131427e-19, 5.7441045e-19, 4.518436e-19, -5.660818e-19, -3.2830325e-19, 8.4127954e-19, 1.3190007e-19, -5.1387163e-19, 2.4095262e-19, 7.3000364e-19, -1.6165998e-19, -2.8164662e-19, 5.852027e-19, 3.7178628e-19, -3.2518403e-19, 1.0274346e-21, 6.2885145e-19, -4.079063e-20, -3.2824618e-19, 2.1637937e-19, 4.2674082e-19, -3.4039816e-19, -2.0769758e-19, 2.9972975e-19, 1.1273107e-19, -4.4162335e-19, -3.7939172e-20, 2.5113276e-19, -1.6912404e-19, -3.5354764e-19, 1.0582358e-19};
	localparam real hb[0:1199] = {0.23903719, 0.056577254, -0.046376806, -0.009240281, 0.16428359, 0.13344508, -0.0036647443, -0.01928589, 0.081619464, 0.15000962, 0.05185026, -0.011636511, 0.014241237, 0.11663765, 0.09115172, 0.010857091, -0.024764504, 0.05822209, 0.098571725, 0.037874848, -0.034566384, 0.0019830666, 0.07477467, 0.058038898, -0.023895573, -0.032810993, 0.03275979, 0.064085096, -0.0055858963, -0.03981509, -0.009921085, 0.055135515, 0.009022917, -0.024662416, -0.03888094, 0.035908896, 0.013744869, 0.00015487392, -0.04764395, 0.013902288, 0.008398102, 0.021689452, -0.03832304, -0.0039017962, -0.0027806722, 0.031541757, -0.018921323, -0.0134365605, -0.013971439, 0.027936192, 0.00094403164, -0.014351925, -0.020490887, 0.01479963, 0.013927031, -0.009275766, -0.020404473, -0.0010919541, 0.017087722, -0.0021609426, -0.014691741, -0.013364744, 0.01189166, 0.003458948, -0.006250252, -0.018378805, 0.0025779814, 0.0056395885, 0.0016081632, -0.015981153, -0.0061094626, 0.004325947, 0.0064796824, -0.008769799, -0.010830792, 0.00087981566, 0.007551678, -0.0004959182, -0.010572402, -0.0028033704, 0.0055375565, 0.0055937036, -0.0064739278, -0.0051599727, 0.0020609503, 0.0078387195, -0.00088632095, -0.005486435, -0.0011527935, 0.0064021344, 0.0038024418, -0.0040134266, -0.0029316158, 0.002772526, 0.0060780346, -0.0016068702, -0.0029507598, -0.0011090921, 0.0056674257, 0.0007025566, -0.001641975, -0.0036829025, 0.003353879, 0.0021434487, 0.00015665147, -0.004262454, 0.00043916042, 0.0024323983, 0.0016177294, -0.0030825865, -0.001862258, 0.0017671462, 0.0022367118, -0.0009908297, -0.0028540406, 0.00064182235, 0.0019474562, 0.0010174464, -0.0024938714, -0.00040492573, 0.0010448572, 0.0022089037, -0.0012531686, -0.0009990553, -1.0437184e-05, 0.0023265942, 0.00018164712, -0.001029527, -0.0008038651, 0.0015748176, 0.0012171555, -0.0006254468, -0.0011118401, 0.00043450092, 0.0015528711, -4.9232138e-05, -0.00094108394, -0.00058160716, 0.0012239799, 0.0004343547, -0.0004725073, -0.001127973, 0.0005082042, 0.0006586299, 4.6858797e-05, -0.0011158069, -0.0002360883, 0.0005945838, 0.00041119408, -0.00068544026, -0.0007235973, 0.00032931016, 0.0005225105, -9.9579425e-05, -0.0008319858, 5.902313e-06, 0.00040127503, 0.0003839079, -0.00060940516, -0.00024349481, 0.00015031172, 0.00060723675, -0.00021633696, -0.00034474264, -0.00010345545, 0.00054791843, 0.00016091713, -0.00029593165, -0.0002623835, 0.0002949932, 0.000385986, -0.000151193, -0.00028780816, -1.084417e-05, 0.00041159766, 1.26556315e-05, -0.00020057078, -0.00024225442, 0.00027615347, 0.00013008782, -5.9104073e-05, -0.00032984538, 6.906533e-05, 0.00016860482, 7.138953e-05, -0.00027448742, -0.00011477901, 0.00013299152, 0.0001450063, -0.0001303883, -0.00021180927, 5.463472e-05, 0.00014781408, 2.7808315e-05, -0.0002061253, -2.6564689e-05, 9.555136e-05, 0.00013779633, -0.0001241317, -7.916516e-05, 2.0756184e-05, 0.00017001014, -1.4608162e-05, -8.995813e-05, -4.3355023e-05, 0.00013094475, 7.487308e-05, -6.459199e-05, -7.5454125e-05, 5.2193198e-05, 0.000115488736, -2.0983176e-05, -7.1249924e-05, -2.7314725e-05, 0.00010352842, 2.030821e-05, -4.1046686e-05, -7.761436e-05, 5.584598e-05, 4.4414155e-05, -2.4226397e-06, -8.679232e-05, -1.3141753e-06, 4.638906e-05, 2.807657e-05, -6.116444e-05, -4.4363027e-05, 3.0722178e-05, 4.088765e-05, -1.8588575e-05, -6.0568334e-05, 7.4315167e-06, 3.535451e-05, 2.095851e-05, -5.0250837e-05, -1.29890805e-05, 1.7861572e-05, 4.3364787e-05, -2.3574563e-05, -2.3606332e-05, -2.2271104e-06, 4.4279313e-05, 5.587432e-06, -2.2796748e-05, -1.6782578e-05, 2.8430753e-05, 2.5723135e-05, -1.3595162e-05, -2.1664937e-05, 5.707431e-06, 3.143047e-05, -1.4546162e-06, -1.7331313e-05, -1.3766452e-05, 2.3991272e-05, 8.367861e-06, -7.57829e-06, -2.3477261e-05, 9.307361e-06, 1.2732551e-05, 2.668597e-06, -2.2106002e-05, -5.4039187e-06, 1.1290444e-05, 9.465061e-06, -1.2792604e-05, -1.46239e-05, 5.9522877e-06, 1.1091634e-05, -9.051408e-07, -1.6196838e-05, -3.626266e-07, 8.170177e-06, 8.496937e-06, -1.1340891e-05, -5.0589033e-06, 2.8765296e-06, 1.2483393e-05, -3.39326e-06, -6.7605965e-06, -2.2419993e-06, 1.08456625e-05, 3.9409356e-06, -5.538049e-06, -5.3080794e-06, 5.5301907e-06, 8.0629225e-06, -2.539449e-06, -5.6583185e-06, -6.0073427e-07, 8.191286e-06, 6.9399124e-07, -3.8039354e-06, -5.0575104e-06, 5.2242754e-06, 2.8979214e-06, -9.610125e-07, -6.567052e-06, 1.0058891e-06, 3.492535e-06, 1.5718692e-06, -5.261336e-06, -2.5883094e-06, 2.6374971e-06, 2.919471e-06, -2.2952581e-06, -4.3607315e-06, 9.970679e-07, 2.857432e-06, 8.2797925e-07, -4.0794885e-06, -6.280356e-07, 1.7422229e-06, 2.9021387e-06, -2.3364687e-06, -1.6326735e-06, 2.402107e-07, 3.399242e-06, -1.3064476e-07, -1.7874688e-06, -9.951585e-07, 2.5066513e-06, 1.6023358e-06, -1.2356509e-06, -1.5649143e-06, 8.875635e-07, 2.3254472e-06, -3.511592e-07, -1.4136614e-06, -6.799244e-07, 2.0069417e-06, 4.560163e-07, -7.6896475e-07, -1.621302e-06, 1.0125854e-06, 9.0188763e-07, 1.0838011e-08, -1.7325017e-06, -1.254113e-07, 9.0496854e-07, 6.017416e-07, -1.1685662e-06, -9.4705706e-07, 5.688418e-07, 8.2722744e-07, -3.0056216e-07, -1.219693e-06, 9.9564744e-08, 6.8940943e-07, 4.7449282e-07, -9.712672e-07, -2.957343e-07, 3.2593118e-07, 8.884072e-07, -4.1816645e-07, -4.8665123e-07, -7.3665895e-08, 8.7171094e-07, 1.6041015e-07, -4.5015815e-07, -3.5119737e-07, 5.326038e-07, 5.418449e-07, -2.5379984e-07, -4.3163485e-07, 7.437376e-08, 6.3004137e-07, -8.962163e-09, -3.3150576e-07, -3.0322713e-07, 4.6143782e-07, 1.8120618e-07, -1.310274e-07, -4.7792867e-07, 1.5998009e-07, 2.58456e-07, 7.100539e-08, -4.32371e-07, -1.3000246e-07, 2.2060979e-07, 1.986052e-07, -2.3576192e-07, -3.026566e-07, 1.0909697e-07, 2.2163921e-07, 2.5306413e-09, -3.2112217e-07, -1.6883664e-08, 1.5625234e-07, 1.8343192e-07, -2.1499358e-07, -1.0673519e-07, 4.786528e-08, 2.528132e-07, -5.3503456e-08, -1.3536831e-07, -5.2761305e-08, 2.1111244e-07, 8.978269e-08, -1.06554204e-07, -1.097939e-07, 1.0024878e-07, 1.6553369e-07, -4.4678764e-08, -1.1220572e-07, -2.189342e-08, 1.613825e-07, 1.9268386e-08, -7.203007e-08, -1.0691534e-07, 9.7803216e-08, 6.085932e-08, -1.439441e-08, -1.3177639e-07, 1.2669572e-08, 6.981926e-08, 3.498757e-08, -1.01415e-07, -5.704394e-08, 5.052182e-08, 5.9581375e-08, -4.027415e-08, -8.889118e-08, 1.6883131e-08, 5.604816e-08, 2.1468104e-08, -7.991713e-08, -1.5107494e-08, 3.2369986e-08, 6.055461e-08, -4.3148642e-08, -3.3864257e-08, 2.18074e-09, 6.771711e-08, 1.0669722e-09, -3.549939e-08, -2.1676367e-08, 4.7833446e-08, 3.441283e-08, -2.345563e-08, -3.1769744e-08, 1.4751694e-08, 4.697896e-08, -5.4814357e-09, -2.7580162e-08, -1.601829e-08, 3.89815e-08, 1.0289445e-08, -1.4058324e-08, -3.3504808e-08, 1.828389e-08, 1.8474266e-08, 1.5237563e-09, -3.4307146e-08, -4.3578865e-09, 1.7804986e-08, 1.2844849e-08, -2.2075891e-08, -2.0006997e-08, 1.0628623e-08, 1.6675804e-08, -4.4765187e-09, -2.4460686e-08, 1.1725421e-09, 1.3356231e-08, 1.0631065e-08, -1.8702641e-08, -6.483426e-09, 5.8222533e-09, 1.8181064e-08, -7.306587e-09, -9.8994235e-09, -2.1075506e-09, 1.7136626e-08, 4.126109e-09, -8.800645e-09, -7.3706787e-09, 9.923937e-09, 1.1306756e-08, -4.6675335e-09, -8.628178e-09, 7.0388245e-10, 1.2554064e-08, 2.3408422e-10, -6.3577685e-09, -6.596456e-09, 8.806126e-09, 3.8872323e-09, -2.2448061e-09, -9.698616e-09, 2.6489575e-09, 5.219948e-09, 1.7346367e-09, -8.435354e-09, -3.0418588e-09, 4.28281e-09, 4.122399e-09, -4.313317e-09, -6.2462773e-09, 1.9641828e-09, 4.401484e-09, 4.473801e-10, -6.3534378e-09, -5.407512e-10, 2.9667435e-09, 3.913248e-09, -4.056658e-09, -2.2500861e-09, 7.611298e-10, 5.093392e-09, -7.850426e-10, -2.7122853e-09, -1.2071054e-09, 4.0872674e-09, 2.0057669e-09, -2.0496311e-09, -2.2573325e-09, 1.7892504e-09, 3.3848249e-09, -7.765635e-10, -2.2137703e-09, -6.344276e-10, 3.170153e-09, 4.85774e-10, -1.3517434e-09, -2.246657e-09, 1.8195114e-09, 1.2673408e-09, -1.8778726e-10, -2.6360196e-09, 1.0753591e-10, 1.3893875e-09, 7.708468e-10, -1.9463269e-09, -1.2392986e-09, 9.623969e-10, 1.2138925e-09, -6.9130207e-10, -1.8032444e-09, 2.7623248e-10, 1.097577e-09, 5.253384e-10, -1.558567e-09, -3.5085534e-10, 5.979019e-10, 1.2572086e-09, -7.883495e-10, -6.980945e-10, -7.28967e-12, 1.3451111e-09, 9.4612825e-11, -7.0175876e-10, -4.664454e-10, 9.086293e-10, 7.3306694e-10, -4.4183632e-10, -6.4225203e-10, 2.3534305e-10, 9.458945e-10, -7.80528e-11, -5.3598964e-10, -3.6661402e-10, 7.5420803e-10, 2.2880702e-10, -2.5423344e-10, -6.8877803e-10, 3.2555897e-10, 3.7734316e-10, 5.5978822e-11, -6.767958e-10, -1.2346603e-10, 3.4943906e-10, 2.7177485e-10, -4.1427922e-10, -4.1994003e-10, 1.9732237e-10, 3.3472522e-10, -5.883345e-11, -4.8899595e-10, 7.354714e-12, 2.5745744e-10, 2.3446747e-10, -3.58634e-10, -1.4038243e-10, 1.0210227e-10, 3.7053643e-10, -1.2488001e-10, -2.0058077e-10, -5.4688632e-11, 3.3566602e-10, 1.002722e-10, -1.71433e-10, -1.5387734e-10, 1.8338935e-10, 2.3456928e-10, -8.500832e-11, -1.7197076e-10, -1.4837351e-12, 2.49249e-10, 1.2775306e-11, -1.213987e-10, -1.420233e-10, 1.6714122e-10, 8.262086e-11, -3.735388e-11, -1.9611368e-10, 4.190402e-11, 1.0499606e-10, 4.0773388e-11, -1.6397626e-10, -6.9364424e-11, 8.2765364e-11, 8.513583e-11, -7.8061155e-11, -1.2831633e-10, 3.481403e-11, 8.712096e-11, 1.6732995e-11, -1.2527049e-10, -1.4815689e-11, 5.6020587e-11, 8.281549e-11, -7.60483e-11, -4.7146446e-11, 1.1312403e-11, 1.0224596e-10, -1.00117145e-11, -5.4170977e-11, -2.7043843e-11, 7.8797455e-11, 4.4135452e-11, -3.9252043e-11, -4.6192872e-11, 3.1402166e-11, 6.893752e-11, -1.3171089e-11, -4.351415e-11, -1.652589e-11, 6.205828e-11, 1.1664765e-11, -2.5179353e-11, -4.691772e-11, 3.3575264e-11, 2.6252545e-11, -1.7598609e-12, -5.2548122e-11, -7.3253437e-13, 2.7557769e-11, 1.6772701e-11, -3.7172775e-11, -2.6641982e-11, 1.8237111e-11, 2.4637521e-11, -1.1521935e-11, -3.6442085e-11, 4.296168e-12, 2.1416377e-11, 1.2368233e-11, -3.0278686e-11, -7.951902e-12, 1.0940336e-11, 2.5970887e-11, -1.4239348e-11, -1.4322662e-11, -1.1507129e-12, 2.662969e-11, 3.332645e-12, -1.38228404e-11, -9.947803e-12, 1.7163118e-11, 1.5495927e-11, -8.2665185e-12, -1.2937575e-11, 3.512875e-12, 1.8977715e-11, -9.312016e-13, -1.0375924e-11, -8.220096e-12, 1.4530316e-11, 5.0157166e-12, -4.536437e-12, -1.4097329e-11, 5.6963457e-12, 7.676661e-12, 1.6185608e-12, -1.33052085e-11, -3.1782758e-12, 6.8335754e-12, 5.7101086e-12, -7.719588e-12, -8.761526e-12, 3.631843e-12, 6.695079e-12, -5.666634e-13, -9.742602e-12, -1.7137145e-13, 4.9403693e-12, 5.104583e-12, -6.8440167e-12, -3.0098257e-12, 1.7516496e-12, 7.5218685e-12, -2.0696214e-12, -4.0493425e-12, -1.3377434e-12, 6.5507734e-12, 2.3489977e-12, -3.326747e-12, -3.194753e-12, 3.3572195e-12, 4.841889e-12, -1.5298277e-12, -3.416e-12, -3.3694139e-13, 4.931802e-12, 4.1430165e-13, -2.3060056e-12, -3.0301805e-12, 3.1541033e-12, 1.7429572e-12, -5.9555876e-13, -3.951248e-12, 6.1656274e-13, 2.1044746e-12, 9.328125e-13, -3.174976e-12, -1.5509085e-12, 1.5925316e-12, 1.7500467e-12, -1.3939086e-12, -2.6245063e-12, 6.056207e-13, 1.7185936e-12, 4.8723834e-13, -2.4613378e-12, -3.7431505e-13, 1.0511981e-12, 1.7405205e-12, -1.4153557e-12, -9.820685e-13, 1.4830509e-13, 2.045425e-12, -8.719608e-14, -1.078248e-12, -5.963031e-13, 1.5123815e-12, 9.590977e-13, -7.479879e-13, -9.413492e-13, 5.3937237e-13, 1.3985704e-12, -2.1590919e-13, -8.522749e-13, -4.0515228e-13, 1.2103922e-12, 2.710028e-13, -4.652271e-13, -9.743356e-13, 6.1363984e-13, 5.4115816e-13, 4.3346716e-15, -1.0439734e-12, -7.152961e-14, 5.447469e-13, 3.6108096e-13, -7.0628827e-13, -5.676717e-13, 3.4354876e-13, 4.9817133e-13, -1.8415388e-13, -7.338075e-13, 6.138003e-14, 4.1629802e-13, 2.8328034e-13, -5.858864e-13, -1.7694975e-13, 1.9796273e-13, 5.339739e-13, -2.5365465e-13, -2.9259809e-13, -4.2781947e-14, 5.25399e-13, 9.4865074e-14, -2.7132075e-13, -2.1050177e-13, 3.2216084e-13, 3.2534034e-13, -1.5350748e-13, -2.5969976e-13, 4.644219e-14, 3.7944105e-13, -6.1238496e-15, -2.0002373e-13, -1.8137262e-13, 2.786792e-13, 1.08651776e-13, -7.959608e-14, -2.8734014e-13, 9.744862e-14, 1.5557243e-13, 4.21126e-14, -2.6064283e-13, -7.7348264e-14, 1.3314051e-13, 1.1923485e-13, -1.426905e-13, -1.8179619e-13, 6.617664e-14, 1.3345648e-13, 7.496745e-16, -1.9345163e-13, -9.704703e-15, 9.4348276e-14, 1.0994244e-13, -1.2992451e-13, -6.398412e-14, 2.9179733e-14, 1.5211905e-13, -3.280078e-14, -8.145635e-14, -3.1480864e-14, 1.2735936e-13, 5.36036e-14, -6.429631e-14, -6.599147e-14, 6.0783206e-14, 9.9479744e-14, -2.7129146e-14, -6.7624685e-14, -1.2783077e-14, 9.725011e-14, 1.1393148e-14, -4.355447e-14, -6.414319e-14, 5.91409e-14, 3.652807e-14, -8.878608e-15, -7.9327875e-14, 7.915383e-15, 4.2035992e-14, 2.0909867e-14, -6.1218805e-14, -3.4143166e-14, 3.0502605e-14, 3.5816368e-14, -2.4479474e-14, -5.346002e-14, 1.0281065e-14, 3.378441e-14, 1.2724337e-14, -4.8188782e-14, -9.000922e-15, 1.958574e-14, 3.6354637e-14, -2.6125325e-14, -2.0347237e-14, 1.4170076e-15, 4.077916e-14, 4.9403117e-16, -2.1389334e-14, -1.2979838e-14, 2.8889444e-14, 2.0624947e-14, -1.4177127e-14, -1.910823e-14, 8.999874e-15, 2.8267477e-14, -3.365282e-15, -1.663186e-14, -9.549115e-15, 2.3517741e-14, 6.1461697e-15, -8.5154204e-15, -2.013078e-14, 1.1088403e-14, 1.1104357e-14, 8.6695934e-16, -2.067033e-14, -2.5488255e-15, 1.07312984e-14, 7.703018e-15, -1.33437556e-14, -1.2002541e-14, 6.429101e-15, 1.0036511e-14, -2.756614e-15, -1.4724213e-14, 7.3880294e-16, 8.060058e-15, 6.3554767e-15, -1.1289081e-14, -3.8806133e-15, 3.5341842e-15, 1.0930514e-14, -4.4410945e-15, -5.953361e-15, -1.2430522e-15, 1.0330117e-14, 2.4478962e-15, -5.306518e-15, -4.4236728e-15, 6.004606e-15, 6.789148e-15, -2.8262453e-15, -5.195027e-15, 4.5543326e-16, 7.560731e-15, 1.2475899e-16, -3.8388605e-15, -3.950191e-15, 5.3190895e-15, 2.3302567e-15, -1.3666794e-15, -5.8337247e-15, 1.6169612e-15, 3.1411114e-15, 1.031731e-15, -5.0872625e-15, -1.8138419e-15, 2.5840159e-15, 2.4759461e-15, -2.613043e-15, -3.7531793e-15, 1.1914624e-15, 2.651249e-15, 2.535249e-16, -3.8282006e-15, -3.1738145e-16, 1.792491e-15, 2.3463746e-15, -2.4522919e-15, -1.3501114e-15, 4.6603213e-16, 3.0652225e-15, -4.841344e-16, -1.6328483e-15, -7.2078856e-16, 2.4663181e-15, 1.1992071e-15, -1.2373428e-15, -1.3567271e-15, 1.0859185e-15, 2.0349842e-15, -4.7226894e-16, -1.3341564e-15, -3.7413691e-16, 1.9110107e-15, 2.884382e-16, -8.174619e-16, -1.348384e-15, 1.1009686e-15, 7.610265e-16, -1.1708761e-16, -1.5871335e-15, 7.057515e-17, 8.367997e-16, 4.612715e-16, -1.1751712e-15, -7.4224137e-16, 5.813567e-16, 7.299883e-16, -4.2081267e-16, -1.084709e-15, 1.6876016e-16, 6.617867e-16, 3.1245285e-16, -9.399971e-16, -2.0931193e-16, 3.61982e-16, 7.551073e-16, -4.7764606e-16, -4.19496e-16, -2.343996e-18, 8.10251e-16, 5.403633e-17, -4.2286145e-16, -2.7951973e-16, 5.4900266e-16, 4.3958625e-16, -2.6712314e-16, -3.8641609e-16, 1.4408786e-16, 5.692695e-16, -4.8260844e-17, -3.2333656e-16, -2.1888496e-16, 4.5512605e-16, 1.3684209e-16, -1.5414671e-16, -4.1396144e-16, 1.9762617e-16, 2.2688286e-16, 3.2686786e-17, -4.0786873e-16, -7.288289e-17, 2.1066367e-16, 1.6304098e-16, -2.5052482e-16, -2.5204995e-16, 1.1941897e-16, 2.0148946e-16, -3.665104e-17, -2.9443006e-16, 5.0741794e-18, 1.5540163e-16, 1.402983e-16, -2.1654863e-16, -8.409328e-17, 6.2049676e-17, 2.2282234e-16, -7.604021e-17, -1.2066377e-16, -3.2426003e-17, 2.0238655e-16, 5.966288e-17, -1.034014e-16, -9.239042e-17, 1.1102243e-16, 1.4089534e-16, -5.1516355e-17, -1.03566977e-16, -2.7007362e-19, 1.5014484e-16, 7.3684595e-18, -7.3324506e-17, -8.51073e-17, 1.0099427e-16, 4.9550762e-17, -2.279296e-17, -1.1799334e-16, 2.5673345e-17, 6.319392e-17, 2.4305675e-17, -9.891874e-17, -4.1422856e-17, 4.9948434e-17, 5.1151986e-17, -4.7328767e-17, -7.7123124e-17, 2.114028e-17, 5.249128e-17, 9.763135e-18, -7.549693e-17, -8.76037e-18, 3.3862246e-17, 4.9680593e-17, -4.5992003e-17, -2.8300896e-17, 6.9675665e-18, 6.154662e-17, -6.2558297e-18, -3.261919e-17, -1.616688e-17, 4.756153e-17, 2.6412777e-17, -2.3703251e-17, -2.7770667e-17, 1.9082496e-17, 4.1457267e-17, -8.02482e-18, -2.6230152e-17, -9.796596e-18, 3.7418835e-17, 6.945198e-18, -1.5234642e-17, -2.8169536e-17, 2.0328207e-17, 1.5770227e-17, -1.1394802e-18, -3.164591e-17, -3.2562355e-19, 1.6601574e-17, 1.0044521e-17, -2.2451783e-17, -1.5966703e-17, 1.1020921e-17, 1.481977e-17, -7.029552e-18, -2.19265e-17, 2.6358658e-18, 1.2916152e-17, 7.372336e-18, -1.826638e-17, -4.7503903e-18, 6.6278893e-18, 1.5603859e-17, -8.634589e-18, -8.609169e-18, -6.525927e-19, 1.6044528e-17, 1.9489192e-18, -8.331167e-18, -5.964738e-18, 1.037425e-17, 9.296625e-18, -5.000055e-18, -7.785942e-18, 2.1628883e-18, 1.1424007e-17, -5.858807e-19, -6.2610566e-18, -4.913737e-18, 8.770813e-18, 3.0023494e-18, -2.753312e-18, -8.4750535e-18, 3.4623657e-18, 4.6168925e-18, 9.545539e-19, -8.020238e-18, -1.8852435e-18, 4.120683e-18, 3.427037e-18, -4.670584e-18, -5.2607545e-18, 2.1993144e-18, 4.0310525e-18, -3.6560315e-19, -5.867471e-18, -9.043013e-20, 2.9829303e-18, 3.056825e-18, -4.133909e-18, -1.8041068e-18, 1.0662837e-18, 4.5244348e-18, -1.2632435e-18, -2.436579e-18, -7.9568426e-19, 3.9506986e-18, 1.4005668e-18, -2.0070983e-18, -1.918856e-18, 2.0337993e-18, 2.9092536e-18, -9.27921e-19, -2.0576966e-18, -1.9057048e-19, 2.9715436e-18, 2.4309225e-19, -1.3933192e-18, -1.8168635e-18, 1.9066255e-18, 1.045802e-18, -3.6464952e-19, -2.377869e-18, 3.8009696e-19, 1.266912e-18, 5.5694417e-19, -1.9158241e-18, -9.272453e-19, 9.613686e-19, 1.0518002e-18, -8.459643e-19, -1.5778744e-18, 3.682704e-19, 1.0357111e-18, 2.8725574e-19, -1.4837246e-18, -2.2225118e-19, 6.3569233e-19, 1.0445882e-18, -8.5640713e-19, -5.897324e-19, 9.2414066e-20, 1.2315208e-18, -5.70255e-20, -6.4941547e-19, -3.568125e-19, 9.131427e-19, 5.7441045e-19, -4.518436e-19, -5.660818e-19, 3.2830325e-19, 8.4127954e-19, -1.3190007e-19, -5.1387163e-19, -2.4095262e-19, 7.3000364e-19, 1.6165998e-19, -2.8164662e-19, -5.852027e-19, 3.7178628e-19, 3.2518403e-19, 1.0274346e-21, -6.2885145e-19, -4.079063e-20, 3.2824618e-19, 2.1637937e-19, -4.2674082e-19, -3.4039816e-19, 2.0769758e-19, 2.9972975e-19, -1.1273107e-19, -4.4162335e-19, 3.7939172e-20, 2.5113276e-19, 1.6912404e-19, -3.5354764e-19, -1.0582358e-19};
endpackage
`endif
