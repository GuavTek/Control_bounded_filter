`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam N = 6;
	localparam M = 6;
	localparam real Lfr[0:5] = {0.9796152, 0.9796152, 0.9612651, 0.9612651, 0.95128894, 0.95128894};
	localparam real Lfi[0:5] = {0.12444234, -0.12444234, 0.087433904, -0.087433904, 0.031214636, -0.031214636};
	localparam real Lbr[0:5] = {0.9796152, 0.9796152, 0.9612651, 0.9612651, 0.95128894, 0.95128894};
	localparam real Lbi[0:5] = {0.12444234, -0.12444234, 0.087433904, -0.087433904, 0.031214636, -0.031214636};
	localparam real Wfr[0:5] = {-9.419306e-06, -9.419306e-06, -6.213538e-06, -6.213538e-06, -2.0324521e-06, -2.0324521e-06};
	localparam real Wfi[0:5] = {6.7119745e-06, -6.7119745e-06, -2.3887221e-06, 2.3887221e-06, -4.975176e-06, 4.975176e-06};
	localparam real Wbr[0:5] = {9.419306e-06, 9.419306e-06, 6.213538e-06, 6.213538e-06, 2.0324521e-06, 2.0324521e-06};
	localparam real Wbi[0:5] = {-6.7119745e-06, 6.7119745e-06, 2.3887221e-06, -2.3887221e-06, 4.975176e-06, -4.975176e-06};
	localparam real Ffr[0:5][0:119] = '{
		'{-402.75336, -14.153609, 19.788008, -0.9162649, -0.44597703, 0.06779118, -406.50742, -0.8980802, 19.298191, -1.2955178, -0.39961275, 0.07261636, -403.70404, 12.04209, 18.513689, -1.6447389, -0.34804708, 0.076166846, -394.55093, 24.468977, 17.4543, -1.9591217, -0.29222926, 0.078417875, -379.3515, 36.19774, 16.143707, -2.2345338, -0.23315269, 0.07936597, -358.49783, 47.05923, 14.608999, -2.4675643, -0.17183778, 0.07902845, -332.46213, 56.90231, 12.880153, -2.6555622, -0.10931518, 0.07744266, -301.78726, 65.59578, 10.989486, -2.7966576, -0.04660913, 0.07466485, -267.07635, 73.03, 8.971088, -2.8897734, 0.015278691, 0.07076885, -228.98175, 79.11806, 6.860231, -2.934622, 0.07538453, 0.06584441, -188.19334, 83.79662, 4.692779, -2.9316907, 0.13279691, 0.059995405, -145.42673, 87.02636, 2.5046055, -2.882214, 0.18666992, 0.053337842, -101.41114, 88.79193, 0.33102107, -2.7881365, 0.23623487, 0.045997694, -56.87756, 89.101685, -1.7937741, -2.6520631, 0.28081077, 0.03810865, -12.547007, 87.986885, -3.8372061, -2.4772022, 0.31981286, 0.02980981, 30.880644, 85.500694, -5.768805, -2.2672985, 0.35275954, 0.021243328, 72.73728, 81.71674, -7.560636, -2.0265613, 0.37927753, 0.01255208, 112.3964, 76.72748, -9.187683, -1.7595857, 0.399105, 0.003877369, 149.28201, 70.64221, -10.628171, -1.4712694, 0.41209307, -0.004643273, 182.87654, 63.584957, -11.863833, -1.1667275, 0.4182053, -0.012878189},
		'{-402.75336, -14.153609, 19.788008, -0.9162649, -0.44597703, 0.06779118, -406.50742, -0.8980802, 19.298191, -1.2955178, -0.39961275, 0.07261636, -403.70404, 12.04209, 18.513689, -1.6447389, -0.34804708, 0.076166846, -394.55093, 24.468977, 17.4543, -1.9591217, -0.29222926, 0.078417875, -379.3515, 36.19774, 16.143707, -2.2345338, -0.23315269, 0.07936597, -358.49783, 47.05923, 14.608999, -2.4675643, -0.17183778, 0.07902845, -332.46213, 56.90231, 12.880153, -2.6555622, -0.10931518, 0.07744266, -301.78726, 65.59578, 10.989486, -2.7966576, -0.04660913, 0.07466485, -267.07635, 73.03, 8.971088, -2.8897734, 0.015278691, 0.07076885, -228.98175, 79.11806, 6.860231, -2.934622, 0.07538453, 0.06584441, -188.19334, 83.79662, 4.692779, -2.9316907, 0.13279691, 0.059995405, -145.42673, 87.02636, 2.5046055, -2.882214, 0.18666992, 0.053337842, -101.41114, 88.79193, 0.33102107, -2.7881365, 0.23623487, 0.045997694, -56.87756, 89.101685, -1.7937741, -2.6520631, 0.28081077, 0.03810865, -12.547007, 87.986885, -3.8372061, -2.4772022, 0.31981286, 0.02980981, 30.880644, 85.500694, -5.768805, -2.2672985, 0.35275954, 0.021243328, 72.73728, 81.71674, -7.560636, -2.0265613, 0.37927753, 0.01255208, 112.3964, 76.72748, -9.187683, -1.7595857, 0.399105, 0.003877369, 149.28201, 70.64221, -10.628171, -1.4712694, 0.41209307, -0.004643273, 182.87654, 63.584957, -11.863833, -1.1667275, 0.4182053, -0.012878189},
		'{-927.919, -79.782906, 30.579605, -6.287539, 0.85779405, 0.0068695024, -962.07776, -57.012863, 28.066689, -6.0978026, 0.9054358, -0.013405413, -985.1044, -35.277195, 25.468796, -5.8652654, 0.94154215, -0.032172456, -997.5488, -14.704, 22.815489, -5.5949774, 0.96657103, -0.049363025, -1000.0203, 4.598006, 20.134819, -5.2919903, 0.9810505, -0.06492762, -993.17773, 22.539158, 17.45317, -4.961309, 0.9855689, -0.078835, -977.7199, 39.048363, 14.795135, -4.60785, 0.9807654, -0.09107122, -954.37695, 54.072475, 12.183405, -4.236402, 0.9673209, -0.10163853, -923.90106, 67.57558, 9.638704, -3.8515904, 0.94594884, -0.11055435, -887.0582, 79.53809, 7.179722, -3.457848, 0.91738623, -0.11784997, -844.6205, 89.955894, 4.82309, -3.059386, 0.88238555, -0.12356937, -797.35815, 98.83924, 2.5833673, -2.6601703, 0.8417068, -0.12776794, -746.0331, 106.21175, 0.47304794, -2.2639034, 0.7961099, -0.1305112, -691.3923, 112.109215, -1.4974104, -1.8740077, 0.74634796, -0.13187349, -634.162, 116.57849, -3.3195438, -1.4936137, 0.6931606, -0.1319367, -575.0424, 119.676285, -4.9868226, -1.1255507, 0.63726825, -0.13078903, -514.7034, 121.46797, -6.4945803, -0.7723424, 0.5793668, -0.12852368, -453.78003, 122.026405, -7.839927, -0.4362038, 0.5201231, -0.12523776, -392.8694, 121.43074, -9.021657, -0.11904267, 0.4601707, -0.121031046, -332.52762, 119.76529, -10.040141, 0.17753714, 0.4001062, -0.116004914},
		'{-927.919, -79.782906, 30.579605, -6.287539, 0.85779405, 0.0068695024, -962.07776, -57.012863, 28.066689, -6.0978026, 0.9054358, -0.013405413, -985.1044, -35.277195, 25.468796, -5.8652654, 0.94154215, -0.032172456, -997.5488, -14.704, 22.815489, -5.5949774, 0.96657103, -0.049363025, -1000.0203, 4.598006, 20.134819, -5.2919903, 0.9810505, -0.06492762, -993.17773, 22.539158, 17.45317, -4.961309, 0.9855689, -0.078835, -977.7199, 39.048363, 14.795135, -4.60785, 0.9807654, -0.09107122, -954.37695, 54.072475, 12.183405, -4.236402, 0.9673209, -0.10163853, -923.90106, 67.57558, 9.638704, -3.8515904, 0.94594884, -0.11055435, -887.0582, 79.53809, 7.179722, -3.457848, 0.91738623, -0.11784997, -844.6205, 89.955894, 4.82309, -3.059386, 0.88238555, -0.12356937, -797.35815, 98.83924, 2.5833673, -2.6601703, 0.8417068, -0.12776794, -746.0331, 106.21175, 0.47304794, -2.2639034, 0.7961099, -0.1305112, -691.3923, 112.109215, -1.4974104, -1.8740077, 0.74634796, -0.13187349, -634.162, 116.57849, -3.3195438, -1.4936137, 0.6931606, -0.1319367, -575.0424, 119.676285, -4.9868226, -1.1255507, 0.63726825, -0.13078903, -514.7034, 121.46797, -6.4945803, -0.7723424, 0.5793668, -0.12852368, -453.78003, 122.026405, -7.839927, -0.4362038, 0.5201231, -0.12523776, -392.8694, 121.43074, -9.021657, -0.11904267, 0.4601707, -0.121031046, -332.52762, 119.76529, -10.040141, 0.17753714, 0.4001062, -0.116004914},
		'{-525.5427, -64.57943, 11.147344, -5.2871203, 1.2039611, -0.29534686, -555.3766, -54.880745, 9.139323, -4.7953863, 1.1078888, -0.2757853, -580.5449, -45.910774, 7.2896175, -4.333862, 1.0171463, -0.2571409, -601.40234, -37.63098, 5.589524, -3.9012494, 0.93153584, -0.2393898, -618.28467, -30.004158, 4.0306573, -3.4962769, 0.85086125, -0.22250736, -631.50934, -22.9944, 2.60495, -3.1176996, 0.77492815, -0.20646839, -641.37616, -16.567118, 1.3046468, -2.7643018, 0.7035447, -0.1912472, -648.16797, -10.689032, 0.12230297, -2.4348972, 0.63652176, -0.17681782, -652.15137, -5.328148, -0.9492213, -2.1283317, 0.57367355, -0.16315405, -653.5772, -0.45375532, -1.9167649, -1.8434824, 0.5148176, -0.1502296, -652.6813, 3.9635978, -2.786871, -1.57926, 0.45977533, -0.13801819, -649.68506, 7.9521217, -3.565794, -1.3346083, 0.40837225, -0.12649359, -644.79614, 11.538809, -4.259505, -1.1085051, 0.36043808, -0.11562979, -638.2089, 14.749456, -4.8736978, -0.8999623, 0.31580687, -0.10540097, -630.1052, 17.608694, -5.4137974, -0.7080259, 0.27431726, -0.09578164, -620.65485, 20.140013, -5.884967, -0.531776, 0.23581265, -0.08674665, -610.0161, 22.365784, -6.2921133, -0.3703269, 0.20014106, -0.07827128, -598.3364, 24.307306, -6.639897, -0.22282659, 0.16715537, -0.070331246, -585.7528, 25.984821, -6.9327383, -0.08845654, 0.13671333, -0.062902756, -572.3924, 27.417547, -7.174826, 0.03356872, 0.10867752, -0.055962566},
		'{-525.5427, -64.57943, 11.147344, -5.2871203, 1.2039611, -0.29534686, -555.3766, -54.880745, 9.139323, -4.7953863, 1.1078888, -0.2757853, -580.5449, -45.910774, 7.2896175, -4.333862, 1.0171463, -0.2571409, -601.40234, -37.63098, 5.589524, -3.9012494, 0.93153584, -0.2393898, -618.28467, -30.004158, 4.0306573, -3.4962769, 0.85086125, -0.22250736, -631.50934, -22.9944, 2.60495, -3.1176996, 0.77492815, -0.20646839, -641.37616, -16.567118, 1.3046468, -2.7643018, 0.7035447, -0.1912472, -648.16797, -10.689032, 0.12230297, -2.4348972, 0.63652176, -0.17681782, -652.15137, -5.328148, -0.9492213, -2.1283317, 0.57367355, -0.16315405, -653.5772, -0.45375532, -1.9167649, -1.8434824, 0.5148176, -0.1502296, -652.6813, 3.9635978, -2.786871, -1.57926, 0.45977533, -0.13801819, -649.68506, 7.9521217, -3.565794, -1.3346083, 0.40837225, -0.12649359, -644.79614, 11.538809, -4.259505, -1.1085051, 0.36043808, -0.11562979, -638.2089, 14.749456, -4.8736978, -0.8999623, 0.31580687, -0.10540097, -630.1052, 17.608694, -5.4137974, -0.7080259, 0.27431726, -0.09578164, -620.65485, 20.140013, -5.884967, -0.531776, 0.23581265, -0.08674665, -610.0161, 22.365784, -6.2921133, -0.3703269, 0.20014106, -0.07827128, -598.3364, 24.307306, -6.639897, -0.22282659, 0.16715537, -0.070331246, -585.7528, 25.984821, -6.9327383, -0.08845654, 0.13671333, -0.062902756, -572.3924, 27.417547, -7.174826, 0.03356872, 0.10867752, -0.055962566}};
	localparam real Ffi[0:5][0:119] = '{
		'{96.1416, -104.20096, 0.6946294, 3.1977122, -0.29952127, -0.049879234, 44.062206, -103.83816, 3.1429353, 3.0185056, -0.348914, -0.040426362, -7.422723, -101.8332, 5.4803796, 2.7957568, -0.39153022, -0.030565731, -57.50929, -98.258804, 7.6725497, 2.5340908, -0.42686075, -0.020464275, -105.435814, -93.210846, 9.688201, 2.2386363, -0.454525, -0.010288612, -150.49393, -86.80624, 11.499669, 1.9149314, -0.47427368, -0.00020239467, -192.03845, -79.18055, 13.083229, 1.5688266, -0.4859896, 0.009636216, -229.49615, -70.48541, 14.419367, 1.206382, -0.48968625, 0.019076928, -262.37305, -60.885693, 15.49299, 0.8337676, -0.48550427, 0.02797952, -290.26022, -50.55653, 16.29355, 0.45716125, -0.47370607, 0.036215805, -312.83835, -39.68031, 16.815115, 0.08265091, -0.45466864, 0.043671384, -329.88043, -28.443588, 17.056322, -0.28386036, -0.42887476, 0.05024712, -341.25314, -17.034008, 17.020311, -0.63674337, -0.39690262, 0.055860333, -346.91663, -5.637297, 16.71455, -0.9707257, -0.35941422, 0.060445692, -346.9228, 5.56564, 16.150606, -1.2809666, -0.3171429, 0.06395585, -341.41223, 16.40148, 15.343869, -1.5631232, -0.27087975, 0.066361725, -330.60974, 26.707045, 14.313204, -1.8134073, -0.22145972, 0.06765253, -314.81876, 36.33165, 13.080569, -2.0286314, -0.16974713, 0.06783546, -294.41437, 45.139183, 11.6705885, -2.2062452, -0.11662131, 0.06693516, -269.8358, 53.009914, 10.110091, -2.3443596, -0.06296218, 0.06499288},
		'{-96.1416, 104.20096, -0.6946294, -3.1977122, 0.29952127, 0.049879234, -44.062206, 103.83816, -3.1429353, -3.0185056, 0.348914, 0.040426362, 7.422723, 101.8332, -5.4803796, -2.7957568, 0.39153022, 0.030565731, 57.50929, 98.258804, -7.6725497, -2.5340908, 0.42686075, 0.020464275, 105.435814, 93.210846, -9.688201, -2.2386363, 0.454525, 0.010288612, 150.49393, 86.80624, -11.499669, -1.9149314, 0.47427368, 0.00020239467, 192.03845, 79.18055, -13.083229, -1.5688266, 0.4859896, -0.009636216, 229.49615, 70.48541, -14.419367, -1.206382, 0.48968625, -0.019076928, 262.37305, 60.885693, -15.49299, -0.8337676, 0.48550427, -0.02797952, 290.26022, 50.55653, -16.29355, -0.45716125, 0.47370607, -0.036215805, 312.83835, 39.68031, -16.815115, -0.08265091, 0.45466864, -0.043671384, 329.88043, 28.443588, -17.056322, 0.28386036, 0.42887476, -0.05024712, 341.25314, 17.034008, -17.020311, 0.63674337, 0.39690262, -0.055860333, 346.91663, 5.637297, -16.71455, 0.9707257, 0.35941422, -0.060445692, 346.9228, -5.56564, -16.150606, 1.2809666, 0.3171429, -0.06395585, 341.41223, -16.40148, -15.343869, 1.5631232, 0.27087975, -0.066361725, 330.60974, -26.707045, -14.313204, 1.8134073, 0.22145972, -0.06765253, 314.81876, -36.33165, -13.080569, 2.0286314, 0.16974713, -0.06783546, 294.41437, -45.139183, -11.6705885, 2.2062452, 0.11662131, -0.06693516, 269.8358, -53.009914, -10.110091, 2.3443596, 0.06296218, -0.06499288},
		'{801.76733, -225.08035, 15.193381, 0.61544776, -0.92490834, 0.22884516, 689.57935, -223.3376, 17.27856, 0.041864358, -0.8140818, 0.22058149, 578.7503, -219.6715, 19.063257, -0.49291196, -0.7033826, 0.2108652, 470.20096, -214.24696, 20.55168, -0.98664206, -0.59381443, 0.19988438, 364.76816, -207.23375, 21.75046, -1.4376153, -0.48630196, 0.18782587, 263.20322, -198.80453, 22.668423, -1.8446287, -0.38168803, 0.17487358, 166.17064, -189.13316, 23.31636, -2.2069638, -0.28073123, 0.161207, 74.24817, -178.39296, 23.7068, -2.5243595, -0.18410498, 0.14699996, -12.072729, -166.75516, 23.853762, -2.7969837, -0.09239704, 0.13241926, -92.38537, -154.38751, 23.772537, -3.0254023, -0.0061100475, 0.11762381, -166.36578, -141.45299, 23.47946, -3.2105467, 0.07433728, 0.102763586, -233.77008, -128.10863, 22.991686, -3.3536804, 0.14860824, 0.08797889, -294.43115, -114.50445, 22.326979, -3.4563649, 0.21644562, 0.07339978, -348.25497, -100.782616, 21.503506, -3.5204248, 0.27766863, 0.059145544, -395.21646, -87.07666, 20.539644, -3.547913, 0.33216926, 0.045324333, -435.35504, -73.51084, 19.453802, -3.5410774, 0.37990844, 0.03203296, -468.76978, -60.19964, 18.264242, -3.5023253, 0.42091155, 0.019356769, -495.61453, -47.24739, 16.988932, -3.434192, 0.45526388, 0.0073696584, -516.0927, -34.74802, 15.645391, -3.3393078, 0.48310566, -0.0038658313, -530.45197, -22.784895, 14.250569, -3.2203681, 0.5046271, -0.014298305},
		'{-801.76733, 225.08035, -15.193381, -0.61544776, 0.92490834, -0.22884516, -689.57935, 223.3376, -17.27856, -0.041864358, 0.8140818, -0.22058149, -578.7503, 219.6715, -19.063257, 0.49291196, 0.7033826, -0.2108652, -470.20096, 214.24696, -20.55168, 0.98664206, 0.59381443, -0.19988438, -364.76816, 207.23375, -21.75046, 1.4376153, 0.48630196, -0.18782587, -263.20322, 198.80453, -22.668423, 1.8446287, 0.38168803, -0.17487358, -166.17064, 189.13316, -23.31636, 2.2069638, 0.28073123, -0.161207, -74.24817, 178.39296, -23.7068, 2.5243595, 0.18410498, -0.14699996, 12.072729, 166.75516, -23.853762, 2.7969837, 0.09239704, -0.13241926, 92.38537, 154.38751, -23.772537, 3.0254023, 0.0061100475, -0.11762381, 166.36578, 141.45299, -23.47946, 3.2105467, -0.07433728, -0.102763586, 233.77008, 128.10863, -22.991686, 3.3536804, -0.14860824, -0.08797889, 294.43115, 114.50445, -22.326979, 3.4563649, -0.21644562, -0.07339978, 348.25497, 100.782616, -21.503506, 3.5204248, -0.27766863, -0.059145544, 395.21646, 87.07666, -20.539644, 3.547913, -0.33216926, -0.045324333, 435.35504, 73.51084, -19.453802, 3.5410774, -0.37990844, -0.03203296, 468.76978, 60.19964, -18.264242, 3.5023253, -0.42091155, -0.019356769, 495.61453, 47.24739, -16.988932, 3.434192, -0.45526388, -0.0073696584, 516.0927, 34.74802, -15.645391, 3.3393078, -0.48310566, 0.0038658313, 530.45197, 22.784895, -14.250569, 3.2203681, -0.5046271, 0.014298305},
		'{1775.8845, -209.93199, 46.93379, -7.502651, 1.1989923, -0.16578464, 1672.9747, -201.72182, 44.995552, -7.3022246, 1.1781694, -0.16692825, 1574.1465, -193.60881, 43.089054, -7.096212, 1.1553618, -0.16740553, 1479.3467, -185.61102, 41.217686, -6.885828, 1.1308328, -0.1672776, 1388.5137, -177.74435, 39.384403, -6.6721883, 1.1048263, -0.16660179, 1301.5781, -170.0228, 37.591763, -6.456314, 1.0775684, -0.16543193, 1218.4646, -162.45857, 35.84194, -6.239138, 1.049268, -0.1638184, 1139.0916, -155.0622, 34.13677, -6.0215096, 1.020118, -0.16180836, 1063.3729, -147.8426, 32.47775, -5.8042, 0.99029577, -0.1594458, 991.21826, -140.80736, 30.866093, -5.587907, 0.9599644, -0.15677182, 922.5338, -133.96265, 29.302742, -5.3732576, 0.9292734, -0.15382467, 857.223, -127.31346, 27.788383, -5.1608167, 0.89835924, -0.1506399, 795.18713, -120.86366, 26.323479, -4.951087, 0.8673464, -0.14725052, 736.3256, -114.61609, 24.908276, -4.7445164, 0.836348, -0.14368714, 680.537, -108.572624, 23.542837, -4.5414977, 0.8054664, -0.13997804, 627.7188, -102.73429, 22.22705, -4.3423777, 0.77479404, -0.13614936, 577.7685, -97.10133, 20.960651, -4.147455, 0.7444138, -0.13222514, 530.5833, -91.67329, 19.743229, -3.9569879, 0.7144, -0.12822753, 486.06122, -86.449036, 18.574255, -3.7711942, 0.6848185, -0.12417679, 444.10062, -81.42691, 17.453081, -3.5902565, 0.65572774, -0.120091505},
		'{-1775.8845, 209.93199, -46.93379, 7.502651, -1.1989923, 0.16578464, -1672.9747, 201.72182, -44.995552, 7.3022246, -1.1781694, 0.16692825, -1574.1465, 193.60881, -43.089054, 7.096212, -1.1553618, 0.16740553, -1479.3467, 185.61102, -41.217686, 6.885828, -1.1308328, 0.1672776, -1388.5137, 177.74435, -39.384403, 6.6721883, -1.1048263, 0.16660179, -1301.5781, 170.0228, -37.591763, 6.456314, -1.0775684, 0.16543193, -1218.4646, 162.45857, -35.84194, 6.239138, -1.049268, 0.1638184, -1139.0916, 155.0622, -34.13677, 6.0215096, -1.020118, 0.16180836, -1063.3729, 147.8426, -32.47775, 5.8042, -0.99029577, 0.1594458, -991.21826, 140.80736, -30.866093, 5.587907, -0.9599644, 0.15677182, -922.5338, 133.96265, -29.302742, 5.3732576, -0.9292734, 0.15382467, -857.223, 127.31346, -27.788383, 5.1608167, -0.89835924, 0.1506399, -795.18713, 120.86366, -26.323479, 4.951087, -0.8673464, 0.14725052, -736.3256, 114.61609, -24.908276, 4.7445164, -0.836348, 0.14368714, -680.537, 108.572624, -23.542837, 4.5414977, -0.8054664, 0.13997804, -627.7188, 102.73429, -22.22705, 4.3423777, -0.77479404, 0.13614936, -577.7685, 97.10133, -20.960651, 4.147455, -0.7444138, 0.13222514, -530.5833, 91.67329, -19.743229, 3.9569879, -0.7144, 0.12822753, -486.06122, 86.449036, -18.574255, 3.7711942, -0.6848185, 0.12417679, -444.10062, 81.42691, -17.453081, 3.5902565, -0.65572774, 0.120091505}};
	localparam real Fbr[0:5][0:119] = '{
		'{402.75336, -14.153609, -19.788008, -0.9162649, 0.44597703, 0.06779118, 406.50742, -0.8980802, -19.298191, -1.2955178, 0.39961275, 0.07261636, 403.70404, 12.04209, -18.513689, -1.6447389, 0.34804708, 0.076166846, 394.55093, 24.468977, -17.4543, -1.9591217, 0.29222926, 0.078417875, 379.3515, 36.19774, -16.143707, -2.2345338, 0.23315269, 0.07936597, 358.49783, 47.05923, -14.608999, -2.4675643, 0.17183778, 0.07902845, 332.46213, 56.90231, -12.880153, -2.6555622, 0.10931518, 0.07744266, 301.78726, 65.59578, -10.989486, -2.7966576, 0.04660913, 0.07466485, 267.07635, 73.03, -8.971088, -2.8897734, -0.015278691, 0.07076885, 228.98175, 79.11806, -6.860231, -2.934622, -0.07538453, 0.06584441, 188.19334, 83.79662, -4.692779, -2.9316907, -0.13279691, 0.059995405, 145.42673, 87.02636, -2.5046055, -2.882214, -0.18666992, 0.053337842, 101.41114, 88.79193, -0.33102107, -2.7881365, -0.23623487, 0.045997694, 56.87756, 89.101685, 1.7937741, -2.6520631, -0.28081077, 0.03810865, 12.547007, 87.986885, 3.8372061, -2.4772022, -0.31981286, 0.02980981, -30.880644, 85.500694, 5.768805, -2.2672985, -0.35275954, 0.021243328, -72.73728, 81.71674, 7.560636, -2.0265613, -0.37927753, 0.01255208, -112.3964, 76.72748, 9.187683, -1.7595857, -0.399105, 0.003877369, -149.28201, 70.64221, 10.628171, -1.4712694, -0.41209307, -0.004643273, -182.87654, 63.584957, 11.863833, -1.1667275, -0.4182053, -0.012878189},
		'{402.75336, -14.153609, -19.788008, -0.9162649, 0.44597703, 0.06779118, 406.50742, -0.8980802, -19.298191, -1.2955178, 0.39961275, 0.07261636, 403.70404, 12.04209, -18.513689, -1.6447389, 0.34804708, 0.076166846, 394.55093, 24.468977, -17.4543, -1.9591217, 0.29222926, 0.078417875, 379.3515, 36.19774, -16.143707, -2.2345338, 0.23315269, 0.07936597, 358.49783, 47.05923, -14.608999, -2.4675643, 0.17183778, 0.07902845, 332.46213, 56.90231, -12.880153, -2.6555622, 0.10931518, 0.07744266, 301.78726, 65.59578, -10.989486, -2.7966576, 0.04660913, 0.07466485, 267.07635, 73.03, -8.971088, -2.8897734, -0.015278691, 0.07076885, 228.98175, 79.11806, -6.860231, -2.934622, -0.07538453, 0.06584441, 188.19334, 83.79662, -4.692779, -2.9316907, -0.13279691, 0.059995405, 145.42673, 87.02636, -2.5046055, -2.882214, -0.18666992, 0.053337842, 101.41114, 88.79193, -0.33102107, -2.7881365, -0.23623487, 0.045997694, 56.87756, 89.101685, 1.7937741, -2.6520631, -0.28081077, 0.03810865, 12.547007, 87.986885, 3.8372061, -2.4772022, -0.31981286, 0.02980981, -30.880644, 85.500694, 5.768805, -2.2672985, -0.35275954, 0.021243328, -72.73728, 81.71674, 7.560636, -2.0265613, -0.37927753, 0.01255208, -112.3964, 76.72748, 9.187683, -1.7595857, -0.399105, 0.003877369, -149.28201, 70.64221, 10.628171, -1.4712694, -0.41209307, -0.004643273, -182.87654, 63.584957, 11.863833, -1.1667275, -0.4182053, -0.012878189},
		'{927.919, -79.782906, -30.579605, -6.287539, -0.85779405, 0.0068695024, 962.07776, -57.012863, -28.066689, -6.0978026, -0.9054358, -0.013405413, 985.1044, -35.277195, -25.468796, -5.8652654, -0.94154215, -0.032172456, 997.5488, -14.704, -22.815489, -5.5949774, -0.96657103, -0.049363025, 1000.0203, 4.598006, -20.134819, -5.2919903, -0.9810505, -0.06492762, 993.17773, 22.539158, -17.45317, -4.961309, -0.9855689, -0.078835, 977.7199, 39.048363, -14.795135, -4.60785, -0.9807654, -0.09107122, 954.37695, 54.072475, -12.183405, -4.236402, -0.9673209, -0.10163853, 923.90106, 67.57558, -9.638704, -3.8515904, -0.94594884, -0.11055435, 887.0582, 79.53809, -7.179722, -3.457848, -0.91738623, -0.11784997, 844.6205, 89.955894, -4.82309, -3.059386, -0.88238555, -0.12356937, 797.35815, 98.83924, -2.5833673, -2.6601703, -0.8417068, -0.12776794, 746.0331, 106.21175, -0.47304794, -2.2639034, -0.7961099, -0.1305112, 691.3923, 112.109215, 1.4974104, -1.8740077, -0.74634796, -0.13187349, 634.162, 116.57849, 3.3195438, -1.4936137, -0.6931606, -0.1319367, 575.0424, 119.676285, 4.9868226, -1.1255507, -0.63726825, -0.13078903, 514.7034, 121.46797, 6.4945803, -0.7723424, -0.5793668, -0.12852368, 453.78003, 122.026405, 7.839927, -0.4362038, -0.5201231, -0.12523776, 392.8694, 121.43074, 9.021657, -0.11904267, -0.4601707, -0.121031046, 332.52762, 119.76529, 10.040141, 0.17753714, -0.4001062, -0.116004914},
		'{927.919, -79.782906, -30.579605, -6.287539, -0.85779405, 0.0068695024, 962.07776, -57.012863, -28.066689, -6.0978026, -0.9054358, -0.013405413, 985.1044, -35.277195, -25.468796, -5.8652654, -0.94154215, -0.032172456, 997.5488, -14.704, -22.815489, -5.5949774, -0.96657103, -0.049363025, 1000.0203, 4.598006, -20.134819, -5.2919903, -0.9810505, -0.06492762, 993.17773, 22.539158, -17.45317, -4.961309, -0.9855689, -0.078835, 977.7199, 39.048363, -14.795135, -4.60785, -0.9807654, -0.09107122, 954.37695, 54.072475, -12.183405, -4.236402, -0.9673209, -0.10163853, 923.90106, 67.57558, -9.638704, -3.8515904, -0.94594884, -0.11055435, 887.0582, 79.53809, -7.179722, -3.457848, -0.91738623, -0.11784997, 844.6205, 89.955894, -4.82309, -3.059386, -0.88238555, -0.12356937, 797.35815, 98.83924, -2.5833673, -2.6601703, -0.8417068, -0.12776794, 746.0331, 106.21175, -0.47304794, -2.2639034, -0.7961099, -0.1305112, 691.3923, 112.109215, 1.4974104, -1.8740077, -0.74634796, -0.13187349, 634.162, 116.57849, 3.3195438, -1.4936137, -0.6931606, -0.1319367, 575.0424, 119.676285, 4.9868226, -1.1255507, -0.63726825, -0.13078903, 514.7034, 121.46797, 6.4945803, -0.7723424, -0.5793668, -0.12852368, 453.78003, 122.026405, 7.839927, -0.4362038, -0.5201231, -0.12523776, 392.8694, 121.43074, 9.021657, -0.11904267, -0.4601707, -0.121031046, 332.52762, 119.76529, 10.040141, 0.17753714, -0.4001062, -0.116004914},
		'{525.5427, -64.57943, -11.147344, -5.2871203, -1.2039611, -0.29534686, 555.3766, -54.880745, -9.139323, -4.7953863, -1.1078888, -0.2757853, 580.5449, -45.910774, -7.2896175, -4.333862, -1.0171463, -0.2571409, 601.40234, -37.63098, -5.589524, -3.9012494, -0.93153584, -0.2393898, 618.28467, -30.004158, -4.0306573, -3.4962769, -0.85086125, -0.22250736, 631.50934, -22.9944, -2.60495, -3.1176996, -0.77492815, -0.20646839, 641.37616, -16.567118, -1.3046468, -2.7643018, -0.7035447, -0.1912472, 648.16797, -10.689032, -0.12230297, -2.4348972, -0.63652176, -0.17681782, 652.15137, -5.328148, 0.9492213, -2.1283317, -0.57367355, -0.16315405, 653.5772, -0.45375532, 1.9167649, -1.8434824, -0.5148176, -0.1502296, 652.6813, 3.9635978, 2.786871, -1.57926, -0.45977533, -0.13801819, 649.68506, 7.9521217, 3.565794, -1.3346083, -0.40837225, -0.12649359, 644.79614, 11.538809, 4.259505, -1.1085051, -0.36043808, -0.11562979, 638.2089, 14.749456, 4.8736978, -0.8999623, -0.31580687, -0.10540097, 630.1052, 17.608694, 5.4137974, -0.7080259, -0.27431726, -0.09578164, 620.65485, 20.140013, 5.884967, -0.531776, -0.23581265, -0.08674665, 610.0161, 22.365784, 6.2921133, -0.3703269, -0.20014106, -0.07827128, 598.3364, 24.307306, 6.639897, -0.22282659, -0.16715537, -0.070331246, 585.7528, 25.984821, 6.9327383, -0.08845654, -0.13671333, -0.062902756, 572.3924, 27.417547, 7.174826, 0.03356872, -0.10867752, -0.055962566},
		'{525.5427, -64.57943, -11.147344, -5.2871203, -1.2039611, -0.29534686, 555.3766, -54.880745, -9.139323, -4.7953863, -1.1078888, -0.2757853, 580.5449, -45.910774, -7.2896175, -4.333862, -1.0171463, -0.2571409, 601.40234, -37.63098, -5.589524, -3.9012494, -0.93153584, -0.2393898, 618.28467, -30.004158, -4.0306573, -3.4962769, -0.85086125, -0.22250736, 631.50934, -22.9944, -2.60495, -3.1176996, -0.77492815, -0.20646839, 641.37616, -16.567118, -1.3046468, -2.7643018, -0.7035447, -0.1912472, 648.16797, -10.689032, -0.12230297, -2.4348972, -0.63652176, -0.17681782, 652.15137, -5.328148, 0.9492213, -2.1283317, -0.57367355, -0.16315405, 653.5772, -0.45375532, 1.9167649, -1.8434824, -0.5148176, -0.1502296, 652.6813, 3.9635978, 2.786871, -1.57926, -0.45977533, -0.13801819, 649.68506, 7.9521217, 3.565794, -1.3346083, -0.40837225, -0.12649359, 644.79614, 11.538809, 4.259505, -1.1085051, -0.36043808, -0.11562979, 638.2089, 14.749456, 4.8736978, -0.8999623, -0.31580687, -0.10540097, 630.1052, 17.608694, 5.4137974, -0.7080259, -0.27431726, -0.09578164, 620.65485, 20.140013, 5.884967, -0.531776, -0.23581265, -0.08674665, 610.0161, 22.365784, 6.2921133, -0.3703269, -0.20014106, -0.07827128, 598.3364, 24.307306, 6.639897, -0.22282659, -0.16715537, -0.070331246, 585.7528, 25.984821, 6.9327383, -0.08845654, -0.13671333, -0.062902756, 572.3924, 27.417547, 7.174826, 0.03356872, -0.10867752, -0.055962566}};
	localparam real Fbi[0:5][0:119] = '{
		'{-96.1416, -104.20096, -0.6946294, 3.1977122, 0.29952127, -0.049879234, -44.062206, -103.83816, -3.1429353, 3.0185056, 0.348914, -0.040426362, 7.422723, -101.8332, -5.4803796, 2.7957568, 0.39153022, -0.030565731, 57.50929, -98.258804, -7.6725497, 2.5340908, 0.42686075, -0.020464275, 105.435814, -93.210846, -9.688201, 2.2386363, 0.454525, -0.010288612, 150.49393, -86.80624, -11.499669, 1.9149314, 0.47427368, -0.00020239467, 192.03845, -79.18055, -13.083229, 1.5688266, 0.4859896, 0.009636216, 229.49615, -70.48541, -14.419367, 1.206382, 0.48968625, 0.019076928, 262.37305, -60.885693, -15.49299, 0.8337676, 0.48550427, 0.02797952, 290.26022, -50.55653, -16.29355, 0.45716125, 0.47370607, 0.036215805, 312.83835, -39.68031, -16.815115, 0.08265091, 0.45466864, 0.043671384, 329.88043, -28.443588, -17.056322, -0.28386036, 0.42887476, 0.05024712, 341.25314, -17.034008, -17.020311, -0.63674337, 0.39690262, 0.055860333, 346.91663, -5.637297, -16.71455, -0.9707257, 0.35941422, 0.060445692, 346.9228, 5.56564, -16.150606, -1.2809666, 0.3171429, 0.06395585, 341.41223, 16.40148, -15.343869, -1.5631232, 0.27087975, 0.066361725, 330.60974, 26.707045, -14.313204, -1.8134073, 0.22145972, 0.06765253, 314.81876, 36.33165, -13.080569, -2.0286314, 0.16974713, 0.06783546, 294.41437, 45.139183, -11.6705885, -2.2062452, 0.11662131, 0.06693516, 269.8358, 53.009914, -10.110091, -2.3443596, 0.06296218, 0.06499288},
		'{96.1416, 104.20096, 0.6946294, -3.1977122, -0.29952127, 0.049879234, 44.062206, 103.83816, 3.1429353, -3.0185056, -0.348914, 0.040426362, -7.422723, 101.8332, 5.4803796, -2.7957568, -0.39153022, 0.030565731, -57.50929, 98.258804, 7.6725497, -2.5340908, -0.42686075, 0.020464275, -105.435814, 93.210846, 9.688201, -2.2386363, -0.454525, 0.010288612, -150.49393, 86.80624, 11.499669, -1.9149314, -0.47427368, 0.00020239467, -192.03845, 79.18055, 13.083229, -1.5688266, -0.4859896, -0.009636216, -229.49615, 70.48541, 14.419367, -1.206382, -0.48968625, -0.019076928, -262.37305, 60.885693, 15.49299, -0.8337676, -0.48550427, -0.02797952, -290.26022, 50.55653, 16.29355, -0.45716125, -0.47370607, -0.036215805, -312.83835, 39.68031, 16.815115, -0.08265091, -0.45466864, -0.043671384, -329.88043, 28.443588, 17.056322, 0.28386036, -0.42887476, -0.05024712, -341.25314, 17.034008, 17.020311, 0.63674337, -0.39690262, -0.055860333, -346.91663, 5.637297, 16.71455, 0.9707257, -0.35941422, -0.060445692, -346.9228, -5.56564, 16.150606, 1.2809666, -0.3171429, -0.06395585, -341.41223, -16.40148, 15.343869, 1.5631232, -0.27087975, -0.066361725, -330.60974, -26.707045, 14.313204, 1.8134073, -0.22145972, -0.06765253, -314.81876, -36.33165, 13.080569, 2.0286314, -0.16974713, -0.06783546, -294.41437, -45.139183, 11.6705885, 2.2062452, -0.11662131, -0.06693516, -269.8358, -53.009914, 10.110091, 2.3443596, -0.06296218, -0.06499288},
		'{-801.76733, -225.08035, -15.193381, 0.61544776, 0.92490834, 0.22884516, -689.57935, -223.3376, -17.27856, 0.041864358, 0.8140818, 0.22058149, -578.7503, -219.6715, -19.063257, -0.49291196, 0.7033826, 0.2108652, -470.20096, -214.24696, -20.55168, -0.98664206, 0.59381443, 0.19988438, -364.76816, -207.23375, -21.75046, -1.4376153, 0.48630196, 0.18782587, -263.20322, -198.80453, -22.668423, -1.8446287, 0.38168803, 0.17487358, -166.17064, -189.13316, -23.31636, -2.2069638, 0.28073123, 0.161207, -74.24817, -178.39296, -23.7068, -2.5243595, 0.18410498, 0.14699996, 12.072729, -166.75516, -23.853762, -2.7969837, 0.09239704, 0.13241926, 92.38537, -154.38751, -23.772537, -3.0254023, 0.0061100475, 0.11762381, 166.36578, -141.45299, -23.47946, -3.2105467, -0.07433728, 0.102763586, 233.77008, -128.10863, -22.991686, -3.3536804, -0.14860824, 0.08797889, 294.43115, -114.50445, -22.326979, -3.4563649, -0.21644562, 0.07339978, 348.25497, -100.782616, -21.503506, -3.5204248, -0.27766863, 0.059145544, 395.21646, -87.07666, -20.539644, -3.547913, -0.33216926, 0.045324333, 435.35504, -73.51084, -19.453802, -3.5410774, -0.37990844, 0.03203296, 468.76978, -60.19964, -18.264242, -3.5023253, -0.42091155, 0.019356769, 495.61453, -47.24739, -16.988932, -3.434192, -0.45526388, 0.0073696584, 516.0927, -34.74802, -15.645391, -3.3393078, -0.48310566, -0.0038658313, 530.45197, -22.784895, -14.250569, -3.2203681, -0.5046271, -0.014298305},
		'{801.76733, 225.08035, 15.193381, -0.61544776, -0.92490834, -0.22884516, 689.57935, 223.3376, 17.27856, -0.041864358, -0.8140818, -0.22058149, 578.7503, 219.6715, 19.063257, 0.49291196, -0.7033826, -0.2108652, 470.20096, 214.24696, 20.55168, 0.98664206, -0.59381443, -0.19988438, 364.76816, 207.23375, 21.75046, 1.4376153, -0.48630196, -0.18782587, 263.20322, 198.80453, 22.668423, 1.8446287, -0.38168803, -0.17487358, 166.17064, 189.13316, 23.31636, 2.2069638, -0.28073123, -0.161207, 74.24817, 178.39296, 23.7068, 2.5243595, -0.18410498, -0.14699996, -12.072729, 166.75516, 23.853762, 2.7969837, -0.09239704, -0.13241926, -92.38537, 154.38751, 23.772537, 3.0254023, -0.0061100475, -0.11762381, -166.36578, 141.45299, 23.47946, 3.2105467, 0.07433728, -0.102763586, -233.77008, 128.10863, 22.991686, 3.3536804, 0.14860824, -0.08797889, -294.43115, 114.50445, 22.326979, 3.4563649, 0.21644562, -0.07339978, -348.25497, 100.782616, 21.503506, 3.5204248, 0.27766863, -0.059145544, -395.21646, 87.07666, 20.539644, 3.547913, 0.33216926, -0.045324333, -435.35504, 73.51084, 19.453802, 3.5410774, 0.37990844, -0.03203296, -468.76978, 60.19964, 18.264242, 3.5023253, 0.42091155, -0.019356769, -495.61453, 47.24739, 16.988932, 3.434192, 0.45526388, -0.0073696584, -516.0927, 34.74802, 15.645391, 3.3393078, 0.48310566, 0.0038658313, -530.45197, 22.784895, 14.250569, 3.2203681, 0.5046271, 0.014298305},
		'{-1775.8845, -209.93199, -46.93379, -7.502651, -1.1989923, -0.16578464, -1672.9747, -201.72182, -44.995552, -7.3022246, -1.1781694, -0.16692825, -1574.1465, -193.60881, -43.089054, -7.096212, -1.1553618, -0.16740553, -1479.3467, -185.61102, -41.217686, -6.885828, -1.1308328, -0.1672776, -1388.5137, -177.74435, -39.384403, -6.6721883, -1.1048263, -0.16660179, -1301.5781, -170.0228, -37.591763, -6.456314, -1.0775684, -0.16543193, -1218.4646, -162.45857, -35.84194, -6.239138, -1.049268, -0.1638184, -1139.0916, -155.0622, -34.13677, -6.0215096, -1.020118, -0.16180836, -1063.3729, -147.8426, -32.47775, -5.8042, -0.99029577, -0.1594458, -991.21826, -140.80736, -30.866093, -5.587907, -0.9599644, -0.15677182, -922.5338, -133.96265, -29.302742, -5.3732576, -0.9292734, -0.15382467, -857.223, -127.31346, -27.788383, -5.1608167, -0.89835924, -0.1506399, -795.18713, -120.86366, -26.323479, -4.951087, -0.8673464, -0.14725052, -736.3256, -114.61609, -24.908276, -4.7445164, -0.836348, -0.14368714, -680.537, -108.572624, -23.542837, -4.5414977, -0.8054664, -0.13997804, -627.7188, -102.73429, -22.22705, -4.3423777, -0.77479404, -0.13614936, -577.7685, -97.10133, -20.960651, -4.147455, -0.7444138, -0.13222514, -530.5833, -91.67329, -19.743229, -3.9569879, -0.7144, -0.12822753, -486.06122, -86.449036, -18.574255, -3.7711942, -0.6848185, -0.12417679, -444.10062, -81.42691, -17.453081, -3.5902565, -0.65572774, -0.120091505},
		'{1775.8845, 209.93199, 46.93379, 7.502651, 1.1989923, 0.16578464, 1672.9747, 201.72182, 44.995552, 7.3022246, 1.1781694, 0.16692825, 1574.1465, 193.60881, 43.089054, 7.096212, 1.1553618, 0.16740553, 1479.3467, 185.61102, 41.217686, 6.885828, 1.1308328, 0.1672776, 1388.5137, 177.74435, 39.384403, 6.6721883, 1.1048263, 0.16660179, 1301.5781, 170.0228, 37.591763, 6.456314, 1.0775684, 0.16543193, 1218.4646, 162.45857, 35.84194, 6.239138, 1.049268, 0.1638184, 1139.0916, 155.0622, 34.13677, 6.0215096, 1.020118, 0.16180836, 1063.3729, 147.8426, 32.47775, 5.8042, 0.99029577, 0.1594458, 991.21826, 140.80736, 30.866093, 5.587907, 0.9599644, 0.15677182, 922.5338, 133.96265, 29.302742, 5.3732576, 0.9292734, 0.15382467, 857.223, 127.31346, 27.788383, 5.1608167, 0.89835924, 0.1506399, 795.18713, 120.86366, 26.323479, 4.951087, 0.8673464, 0.14725052, 736.3256, 114.61609, 24.908276, 4.7445164, 0.836348, 0.14368714, 680.537, 108.572624, 23.542837, 4.5414977, 0.8054664, 0.13997804, 627.7188, 102.73429, 22.22705, 4.3423777, 0.77479404, 0.13614936, 577.7685, 97.10133, 20.960651, 4.147455, 0.7444138, 0.13222514, 530.5833, 91.67329, 19.743229, 3.9569879, 0.7144, 0.12822753, 486.06122, 86.449036, 18.574255, 3.7711942, 0.6848185, 0.12417679, 444.10062, 81.42691, 17.453081, 3.5902565, 0.65572774, 0.120091505}};
	localparam real hf[0:1799] = {0.04146539, -0.00024480597, -0.00026783795, 2.248845e-06, 4.3801842e-06, -4.864713e-08, 0.041221026, -0.00073176116, -0.0002614101, 6.696438e-06, 4.290541e-06, -1.448581e-07, 0.040734954, -0.0012107815, -0.00024864986, 1.0994666e-05, 4.1132726e-06, -2.3784936e-07, 0.04001243, -0.0016766941, -0.0002297464, 1.5047003e-05, 3.8523635e-06, -3.2557224e-07, 0.039061278, -0.0021244998, -0.00020497982, 1.8761422e-05, 3.5136645e-06, -4.06118e-07, 0.037891746, -0.0025494383, -0.00017471658, 2.205205e-05, 3.1047541e-06, -4.7776365e-07, 0.036516394, -0.0029470513, -0.00013940375, 2.4840714e-05, 2.6347661e-06, -5.3901107e-07, 0.034949932, -0.0033132397, -9.9561985e-05, 2.7058317e-05, 2.1141852e-06, -5.8861855e-07, 0.03320901, -0.003644315, -5.5777306e-05, 2.8646065e-05, 1.5546185e-06, -6.256258e-07, 0.03131201, -0.003937048, -8.692036e-06, 2.9556486e-05, 9.685473e-07, -6.493704e-07, 0.029278811, -0.0041887052, 4.100521e-05, 2.9754228e-05, 3.690637e-07, -6.594982e-07, 0.027130522, -0.0043970835, 9.259013e-05, 2.9216664e-05, -2.3039931e-07, -6.559652e-07, 0.024889218, -0.0045605334, 0.00014531388, 2.7934244e-05, -8.163425e-07, -6.390335e-07, 0.02257766, -0.004677976, 0.00019841442, 2.5910616e-05, -1.3754711e-06, -6.092603e-07, 0.020218996, -0.0047489107, 0.00025112805, 2.3162525e-05, -1.8949582e-06, -5.6748127e-07, 0.01783649, -0.0047734166, 0.00030270085, 1.9719477e-05, -2.3626956e-06, -5.1478764e-07, 0.015453213, -0.0047521433, 0.00035239992, 1.5623187e-05, -2.7675267e-06, -4.5249982e-07, 0.013091778, -0.004686295, 0.00039952397, 1.0926819e-05, -3.0994586e-06, -3.8213585e-07, 0.010774061, -0.0045776074, 0.00044341368, 5.6940457e-06, -3.34985e-06, -3.053772e-07, 0.008520941, -0.004428317, 0.00048346096, -2.079197e-09, -3.5115697e-06, -2.2403161e-07, 0.0063520637, -0.004241123, 0.0005191175, -6.08038e-06, -3.579126e-06, -1.3999463e-07, 0.0042856177, -0.004019145, 0.0005499023, -1.2452956e-05, -3.548764e-06, -5.5209913e-08, 0.0023381365, -0.0037658734, 0.000575408, -1.902667e-05, -3.4185289e-06, 2.8370449e-08, 0.00052432675, -0.0034851169, 0.00059530616, -2.5704714e-05, -3.1882964e-06, 1.0882508e-07, -0.0011430768, -0.0031809455, 0.0006093511, -3.2388223e-05, -2.8597694e-06, 1.8430102e-07, -0.0026534274, -0.0028576308, 0.0006173824, -3.8977894e-05, -2.4364408e-06, 2.5304948e-07, -0.0039982516, -0.002519585, 0.0006193266, -4.5375622e-05, -1.9235256e-06, 3.1345897e-07, -0.0051713055, -0.0021712987, 0.00061519654, -5.1486055e-05, -1.3278617e-06, 3.640851e-07, -0.006168595, -0.0018172781, 0.0006050904, -5.721813e-05, -6.577848e-07, 4.036769e-07, -0.0069883717, -0.0014619845, 0.0005891891, -6.248652e-05, 7.702353e-08, 4.3119886e-07, -0.007631094, -0.001109774, 0.0005677523, -6.721291e-05, 8.65709e-07, 4.4584894e-07, -0.00809936, -0.0007648413, 0.00054111326, -7.132724e-05, 1.6964362e-06, 4.4707144e-07, -0.008397813, -0.00043116606, 0.00050967326, -7.476873e-05, 2.5565953e-06, 4.345657e-07, -0.008533023, -0.000112463655, 0.00047389444, -7.748676e-05, 3.43302e-06, 4.0828954e-07, -0.008513342, 0.00018785929, 0.00043429201, -7.9441576e-05, 4.3122127e-06, 3.684583e-07, -0.008348739, 0.00046674386, 0.00039142597, -8.0604856e-05, 5.180572e-06, 3.1553893e-07, -0.00805062, 0.00072151225, 0.00034589216, -8.096e-05, 6.0246216e-06, 2.5023982e-07, -0.007631627, 0.0009498948, 0.000298313, -8.05023e-05, 6.831232e-06, 1.7349653e-07, -0.007105432, 0.0011500503, 0.00024932786, -7.923891e-05, 7.5878356e-06, 8.645332e-08, -0.0064865164, 0.0013205807, 0.00019958348, -7.71886e-05, 8.282629e-06, -9.558333e-09, -0.0057899496, 0.0014605374, 0.00014972452, -7.4381336e-05, 8.904762e-06, -1.1304449e-07, -0.00503116, 0.001569423, 0.00010038412, -7.085774e-05, 9.444505e-06, -2.2237596e-07, -0.004225716, 0.0016471844, 5.217493e-05, -6.6668326e-05, 9.893401e-06, -3.3581745e-07, -0.0033891022, 0.0016942013, 5.6806734e-06, -6.187262e-05, 1.0244392e-05, -4.5155824e-07, -0.0025365087, 0.0017112679, -3.8551792e-05, -5.6538138e-05, 1.0491919e-05, -5.6774377e-07, -0.0016826305, 0.0016995692, -8.001964e-05, -5.07393e-05, 1.0632002e-05, -6.825074e-07, -0.0008414778, 0.0016606523, -0.00011827045, -4.4556207e-05, 1.06622865e-05, -7.9400235e-07, -2.6203514e-05, 0.0015963936, -0.0001529077, -3.807334e-05, 1.0582069e-05, -9.0043227e-07, 0.00075105205, 0.0015089608, -0.00018359527, -3.1378277e-05, 1.0392294e-05, -1.0000812e-06, 0.0014792971, 0.0014007733, -0.00021006101, -2.4560304e-05, 1.009552e-05, -1.0913416e-06, 0.002148803, 0.0012744586, -0.00023209922, -1.7709088e-05, 9.695872e-06, -1.1727395e-06, 0.0027511988, 0.0011328079, -0.00024957207, -1.0913319e-05, 9.1989505e-06, -1.2429585e-06, 0.0032795395, 0.0009787299, -0.00026241003, -4.2594206e-06, 8.61174e-06, -1.3008598e-06, 0.0037283541, 0.0008152043, -0.00027061123, 2.169698e-06, 7.942478e-06, -1.3454986e-06, 0.00409367, 0.0006452354, -0.00027423972, 8.295808e-06, 7.2005223e-06, -1.3761386e-06, 0.0043730135, 0.0004718075, -0.00027342307, 1.4046433e-05, 6.396189e-06, -1.3922617e-06, 0.004565388, 0.00029784048, -0.00026834864, 1.935582e-05, 5.5405853e-06, -1.393574e-06, 0.0046712337, 0.00012614891, -0.00025925948, 2.4165789e-05, 4.645431e-06, -1.3800093e-06, 0.004692362, -4.059674e-05, -0.0002464492, 2.8426433e-05, 3.7228735e-06, -1.3517264e-06, 0.004631878, -0.00019990538, -0.00023025631, 3.2096712e-05, 2.785297e-06, -1.3091061e-06, 0.004494078, -0.0003494969, -0.00021105794, 3.514487e-05, 1.8451333e-06, -1.2527415e-06, 0.0042843423, -0.0004873296, -0.0001892633, 3.7548714e-05, 9.1467405e-07, -1.1834273e-06, 0.004009006, -0.0006116232, -0.00016530664, 3.929575e-05, 5.888459e-09, -1.1021446e-06, 0.003675227, -0.0007208773, -0.00013964009, 4.038316e-05, -8.697514e-07, -1.0100435e-06, 0.0032908383, -0.0008138848, -0.00011272643, 4.0817617e-05, -1.701434e-06, -9.08424e-07, 0.0028642027, -0.0008897404, -8.5031825e-05, 4.0615e-05, -2.4791593e-06, -7.9871296e-07, 0.0024040581, -0.00094784505, -5.701874e-05, 3.9799936e-05, -3.1938737e-06, -6.8244145e-07, 0.0019193669, -0.0009879041, -2.9139079e-05, 3.8405236e-05, -3.837589e-06, -5.6121934e-07, 0.0014191625, -0.0010099224, -1.8276651e-06, 3.647122e-05, -4.4034823e-06, -4.367096e-07, 0.0009124039, -0.0010141934, 2.450384e-05, 3.4044948e-05, -4.885976e-06, -3.1060247e-07, 0.00040783366, -0.0010012859, 4.9472517e-05, 3.1179337e-05, -5.2807973e-06, -1.845891e-07, -8.6154956e-05, -0.00097202475, 7.272916e-05, 2.793225e-05, -5.585017e-06, -6.033577e-08, -0.000561641, -0.0009274706, 9.396263e-05, 2.4365498e-05, -5.797066e-06, 6.0540856e-08, -0.0010112876, -0.0008688947, 0.000112903464, 2.0543823e-05, -5.916733e-06, 1.7649754e-07, -0.0014284403, -0.0007977517, 0.00012932679, 1.6533855e-05, -5.9451363e-06, 2.8608656e-07, -0.0018072124, -0.00071565114, 0.00014305445, 1.240306e-05, -5.884684e-06, 3.8797606e-07, -0.0021425537, -0.0006243265, 0.00015395635, 8.218712e-06, -5.7390066e-06, 4.809681e-07, -0.0024303054, -0.00052560354, 0.00016195106, 4.046875e-06, -5.5128776e-06, 5.640142e-07, -0.0026672382, -0.00042136834, 0.00016700556, -4.855194e-08, -5.212119e-06, 6.36229e-07, -0.002851074, -0.0003135352, 0.00016913444, -4.006748e-06, -4.8434886e-06, 6.9689986e-07, -0.0029804923, -0.00020401487, 0.00016839804, -7.770807e-06, -4.4145577e-06, 7.454949e-07, -0.0030551208, -9.468427e-05, 0.00016490035, -1.1288498e-05, -3.9335814e-06, 7.816673e-07, -0.0030755112, 1.2642788e-05, 0.00015878597, -1.451293e-05, -3.4093562e-06, 8.05257e-07, -0.0030431, 0.000116242794, 0.00015023665, -1.7403117e-05, -2.8510776e-06, 8.162893e-07, -0.0029601583, 0.00021450751, 0.00013946736, -1.9924453e-05, -2.2681913e-06, 8.1497086e-07, -0.0028297275, 0.0003059664, 0.00012672189, -2.2049056e-05, -1.6702459e-06, 8.0168275e-07, -0.002655546, 0.0003893061, 0.0001122682, -2.3756009e-05, -1.066746e-06, 7.769712e-07, -0.0024419657, 0.00046338706, 9.639343e-05, -2.5031492e-05, -4.6701115e-07, 7.415358e-07, -0.002193862, 0.0005272565, 7.939882e-05, -2.58688e-05, 1.1996097e-07, 6.9621575e-07, -0.0019165382, 0.00058015855, 6.159456e-05, -2.6268237e-05, 6.856217e-07, 6.4197405e-07, -0.0016156246, 0.00062154036, 4.3294538e-05, -2.6236929e-05, 1.2219896e-06, 5.798804e-07, -0.0012969768, 0.00065105513, 2.4811325e-05, -2.578851e-05, 1.7217562e-06, 5.1109276e-07, -0.00096657197, 0.0006685619, 6.4511933e-06, -2.4942734e-05, 2.1783806e-06, 4.368377e-07, -0.0006304072, 0.0006741216, -1.1490546e-05, -2.3725e-05, 2.5861673e-06, 3.5839042e-07, -0.00029439994, 0.0006679901, -2.8733944e-05, -2.2165796e-05, 2.9403316e-06, 2.770545e-07, 3.570702e-05, 0.00065060885, -4.5018438e-05, -2.030007e-05, 3.2370483e-06, 1.9414136e-07, 0.0003544354, 0.00062259194, -6.0106442e-05, -1.8166582e-05, 3.4734844e-06, 1.10950424e-07, 0.0006566542, 0.00058471126, -7.378651e-05, -1.580717e-05, 3.6478157e-06, 2.8749648e-08, 0.0009376542, 0.0005378797, -8.587597e-05, -1.32660225e-05, 3.759228e-06, -5.124282e-08, 0.001193214, 0.0004831321, -9.6223e-05, -1.0588912e-05, 3.8079017e-06, -1.2787592e-07, 0.0014196559, 0.00042160501, -0.00010470825, -7.822441e-06, 3.794983e-06, -2.0008146e-07, 0.0016138916, 0.0003545153, -0.000111245805, -5.0132785e-06, 3.7225384e-06, -2.668882e-07, 0.0017734565, 0.0002831382, -0.000115783645, -2.2074303e-06, 3.5934993e-06, -3.2743432e-07, 0.0018965335, 0.00020878478, -0.00011830353, 5.504701e-07, 3.411592e-06, -3.8097758e-07, 0.001981966, 0.00013277972, -0.000118820346, 3.2178243e-06, 3.1812583e-06, -4.269036e-07, 0.0020292576, 5.6439232e-05, -0.000117380994, 5.7546863e-06, 2.907567e-06, -4.6473204e-07, 0.002038564, -1.895013e-05, -0.00011406272, 8.124317e-06, 2.5961187e-06, -4.941203e-07, 0.0020106724, -9.2151655e-05, -0.00010897106, 1.0293679e-05, 2.2529423e-06, -5.148652e-07, 0.0019469721, -0.0001619973, -0.00010223735, 1.2233855e-05, 1.8843914e-06, -5.269025e-07, 0.0018494154, -0.00022740495, -9.401595e-05, 1.3920389e-05, 1.4970343e-06, -5.3030413e-07, 0.001720471, -0.00028739372, -8.448112e-05, 1.5333557e-05, 1.097547e-06, -5.252735e-07, 0.0015630699, -0.0003410973, -7.382368e-05, 1.6458544e-05, 6.926051e-07, -5.121386e-07, 0.0013805453, -0.00038777513, -6.22475e-05, 1.7285545e-05, 2.887793e-07, -4.9134405e-07, 0.0011765675, -0.00042682106, -4.9965845e-05, 1.7809787e-05, -1.0756439e-07, -4.6344078e-07, 0.0009550746, -0.0004577699, -3.719775e-05, 1.803146e-05, -4.90359e-07, -4.2907462e-07, 0.00072020135, -0.00048030124, -2.4164285e-05, 1.7955588e-05, -8.539238e-07, -3.8897377e-07, 0.00047620616, -0.0004942409, -1.10849605e-05, 1.7591809e-05, -1.1930427e-06, -3.4393543e-07, 0.000227398, -0.0004995602, 1.8257559e-06, 1.6954098e-05, -1.503034e-06, -2.9481123e-07, -2.1935415e-05, -0.0004963725, 1.4361768e-05, 1.6060432e-05, -1.7798089e-06, -2.4249272e-07, -0.0002675976, -0.00048492796, 2.6328446e-05, 1.4932386e-05, -2.0199202e-06, -1.8789628e-07, -0.0005055498, -0.00046560587, 3.7545466e-05, 1.35947e-05, -2.2205988e-06, -1.3194817e-07, -0.0007319731, -0.00043890523, 4.7849324e-05, 1.2074796e-05, -2.379779e-06, -7.556981e-08, -0.000943326, -0.0004054338, 5.7095556e-05, 1.0402267e-05, -2.496112e-06, -1.966345e-08, -0.0011363953, -0.00036589528, 6.516055e-05, 8.608349e-06, -2.5689671e-06, 3.490142e-08, -0.0013083407, -0.00032107567, 7.194299e-05, 6.7253745e-06, -2.5984232e-06, 8.7300805e-08, -0.0014567326, -0.0002718284, 7.736494e-05, 4.7862313e-06, -2.585247e-06, 1.3676791e-07, -0.0015795819, -0.00021905889, 8.1372455e-05, 2.823819e-06, -2.5308632e-06, 1.8260363e-07, -0.0016753613, -0.00016370844, 8.393588e-05, 8.705237e-07, -2.4373128e-06, 2.2418568e-07, -0.0017430203, -0.00010673826, 8.504967e-05, -1.0422855e-06, -2.3072055e-06, 2.6097635e-07, -0.0017819905, -4.9113318e-05, 8.473187e-05, -2.884732e-06, -2.1436617e-06, 2.9252863e-07, -0.0017921835, 8.213343e-06, 8.302324e-05, -4.62887e-06, -1.9502497e-06, 3.184908e-07, -0.0017739814, 6.431576e-05, 7.998597e-05, -6.249081e-06, -1.7309167e-06, 3.386095e-07, -0.0017282194, 0.00011830935, 7.5702206e-05, -7.7224195e-06, -1.4899155e-06, 3.527309e-07, -0.0016561622, 0.00016936421, 7.027217e-05, -9.028916e-06, -1.2317291e-06, 3.6080053e-07, -0.0015594726, 0.00021671722, 6.381213e-05, -1.0151813e-05, -9.609931e-07, 3.6286144e-07, -0.0014401767, 0.00025968274, 5.6452052e-05, -1.1077749e-05, -6.824175e-07, 3.5905097e-07, -0.0013006215, 0.00029766184, 4.8333266e-05, -1.1796891e-05, -4.0070975e-07, 3.4959587e-07, -0.0011434306, 0.00033014987, 3.9605828e-05, -1.230299e-05, -1.2049978e-07, 3.3480643e-07, -0.00097145484, 0.0003567423, 3.0425923e-05, -1.2593396e-05, 1.537317e-07, 3.150693e-07, -0.00078772154, 0.00037713893, 2.0953192e-05, -1.2668999e-05, 4.1772083e-07, 2.9083918e-07, -0.0005953814, 0.0003911462, 1.134808e-05, -1.2534132e-05, 6.6748277e-07, 2.6263004e-07, -0.00039765524, 0.00039867766, 1.7692399e-06, -1.2196404e-05, 8.99368e-07, 2.3100505e-07, -0.00019778035, 0.00039975307, -7.628977e-06, -1.1666498e-05, 1.1101118e-06, 1.965666e-07, 1.0417496e-06, 0.00039449532, -1.669889e-05, -1.0957918e-05, 1.296876e-06, 1.599455e-07, 0.00019569589, 0.0003831261, -2.5301697e-05, -1.0086704e-05, 1.4572834e-06, 1.2179028e-07, 0.00038320126, 0.00036596006, -3.3309487e-05, -9.071102e-06, 1.5894433e-06, 8.275637e-08, 0.0005607561, 0.00034339743, -4.0607014e-05, -7.931223e-06, 1.6919691e-06, 4.349549e-08, 0.00072577846, 0.00031591573, -4.709325e-05, -6.6886664e-06, 1.7639875e-06, 4.645376e-09, 0.0008759425, 0.0002840602, -5.2682648e-05, -5.3661397e-06, 1.8051384e-06, -3.3179994e-08, 0.0010092098, 0.0002484334, -5.7306126e-05, -3.987063e-06, 1.8155679e-06, -6.939956e-08, 0.0011238554, 0.00020968445, -6.091179e-05, -2.5751765e-06, 1.7959125e-06, -1.0347359e-07, 0.0012184877, 0.00016849731, -6.346532e-05, -1.1541526e-06, 1.7472757e-06, -1.3491113e-07, 0.0012920641, 0.00012557908, -6.4950116e-05, 2.5278408e-07, 1.6711991e-06, -1.6327662e-07, 0.0013438981, 8.164823e-05, -6.5367116e-05, 1.623217e-06, 1.5696256e-06, -1.8819536e-07, 0.0013736633, 3.742277e-05, -6.473434e-05, 2.9358766e-06, 1.4448581e-06, -2.0935782e-07, 0.0013813896, -6.3911475e-06, -6.308622e-05, 4.170953e-06, 1.2995133e-06, -2.26523e-07, 0.0013674548, -4.9110262e-05, -6.047262e-05, 5.310377e-06, 1.136472e-06, -2.3952038e-07, 0.0013325703, -9.008453e-05, -5.695766e-05, 6.3380653e-06, 9.588255e-07, -2.4825076e-07, 0.0012777626, -0.00012870673, -5.261836e-05, 7.24013e-06, 7.6982104e-07, -2.5268616e-07, 0.0012043486, -0.00016442109, -4.7543097e-05, 8.005044e-06, 5.7280613e-07, -2.528682e-07, 0.0011139092, -0.00019673095, -4.182989e-05, 8.623769e-06, 3.7117152e-07, -2.4890576e-07, 0.0010082573, -0.00022520528, -3.558463e-05, 9.089839e-06, 1.6829631e-07, -2.4097142e-07, 0.00088940363, -0.00024948397, -2.8919168e-05, 9.399396e-06, -3.250605e-08, -2.2929709e-07, 0.00075952057, -0.00026928185, -2.1949405e-05, 9.5511905e-06, -2.2803921e-07, -2.1416871e-07, 0.0006209036, -0.00028439148, -1.4793331e-05, 9.546537e-06, -4.1527218e-07, -1.9592031e-07, 0.00047593226, -0.00029468464, -7.569097e-06, 9.389224e-06, -5.9138364e-07, -1.7492742e-07, 0.0003270303, -0.00030011236, -3.9312047e-07, 9.0854e-06, -7.5380206e-07, -1.5160002e-07, 0.00017662637, -0.0003007039, 6.621728e-06, 8.643411e-06, -9.002402e-07, -1.2637503e-07, 2.7115331e-05, -0.00029656442, 1.3367841e-05, 8.073614e-06, -1.0287251e-06, -9.970865e-08, -0.000119178745, -0.00028787146, 1.9744464e-05, 7.3881624e-06, -1.1376214e-06, -7.206857e-08, -0.00026003775, -0.0002748704, 2.565913e-05, 6.6007674e-06, -1.2256492e-06, -4.392621e-08, -0.0003933821, -0.00025786896, 3.1028943e-05, 5.7264383e-06, -1.2918955e-06, -1.5749015e-08, -0.00051730033, -0.0002372308, 3.5781653e-05, 4.7812127e-06, -1.3358201e-06, 1.2006875e-08, -0.0006300753, -0.00021336837, 3.9856568e-05, 3.781874e-06, -1.3572542e-06, 3.890365e-08, -0.0007302067, -0.0001867353, 4.320522e-05, 2.7456647e-06, -1.3563944e-06, 6.452839e-08, -0.00081642973, -0.00015781808, 4.5791854e-05, 1.6899994e-06, -1.3337901e-06, 8.849904e-08, -0.00088772917, -0.00012712766, 4.759369e-05, 6.3218243e-07, -1.2903263e-06, 1.10469735e-07, -0.0009433496, -9.51907e-05, 4.8600963e-05, -4.108655e-07, -1.2272005e-06, 1.3013542e-07, -0.0009828011, -6.254085e-05, 4.881676e-05, -1.4228688e-06, -1.1458965e-06, 1.4723571e-07, -0.0010058604, -2.9710145e-05, 4.8256672e-05, -2.3884404e-06, -1.0481527e-06, 1.6155796e-07, -0.0010125681, 2.7794342e-06, 4.6948237e-05, -3.2933067e-06, -9.359288e-07, 1.7293941e-07, -0.001003222, 3.4423952e-05, 4.49302e-05, -4.124507e-06, -8.1136835e-07, 1.8126859e-07, -0.000978365, 6.474508e-05, 4.225164e-05, -4.870569e-06, -6.767601e-07, 1.8648575e-07, -0.00093877193, 9.3297065e-05, 3.8970928e-05, -5.521654e-06, -5.344981e-07, 1.885826e-07, -0.00088543084, 0.000119672986, 3.5154586e-05, -6.0696775e-06, -3.870403e-07, 1.8760112e-07, -0.0008195223, 0.00014351026, 3.0876014e-05, -6.508391e-06, -2.3686813e-07, 1.8363157e-07, -0.0007423962, 0.0001644953, 2.6214162e-05, -6.833439e-06, -8.644602e-08, 1.7680995e-07, -0.00065554614, 0.00018236731, 2.1252148e-05, -7.0423816e-06, 6.181753e-08, 1.6731461e-07, -0.00056058227, 0.00019692112, 1.6075826e-05, -7.134687e-06, 2.0560704e-07, 1.5536234e-07, -0.000459203, 0.00020800902, 1.0772361e-05, -7.111694e-06, 3.427347e-07, 1.4120398e-07, -0.0003531661, 0.00021554178, 5.4288053e-06, -6.976542e-06, 4.7117229e-07, 1.2511956e-07, -0.00024425922, 0.00021948859, 1.3072744e-07, -6.734081e-06, 5.890795e-07, 1.0741304e-07, -0.00013427105, 0.00021987609, -5.0391163e-06, -6.39075e-06, 6.948289e-07, 8.840692e-08, -2.4962921e-05, 0.0002167866, -1.0002027e-05, -5.954436e-06, 7.870264e-07, 6.843662e-08, 8.195832e-05, 0.00021035537, -1.46845105e-05, -5.434313e-06, 8.645281e-07, 4.7844743e-08, 0.00018486603, 0.0002007672, -1.901932e-05, -4.8406664e-06, 9.264522e-07, 2.6975489e-08, 0.00028223748, 0.00018825223, -2.2946373e-05, -4.184698e-06, 9.721866e-07, 6.1690666e-09, 0.0003726754, 0.00017308127, -2.641352e-05, -3.4783302e-06, 1.0013924e-06, -1.4243616e-08, 0.00045492692, 0.00015556037, -2.9377186e-05, -2.7339945e-06, 1.0140021e-06, -3.394602e-08, 0.00052789995, 0.00013602525, -3.1802854e-05, -1.964424e-06, 1.0102143e-06, -5.2640676e-08, 0.00059067627, 0.00011483514, -3.3665376e-05, -1.1824418e-06, 9.904842e-07, -7.005346e-08, 0.00064252195, 9.236654e-05, -3.4949164e-05, -4.0075614e-07, 9.555097e-07, -8.5937394e-08, 0.00068289426, 6.900684e-05, -3.564818e-05, 3.6824008e-07, 9.0621444e-07, -1.0007594e-07, 0.0007114456, 4.5147888e-05, -3.5765814e-05, 1.112658e-06, 8.4372783e-07, -1.1228567e-07, 0.00072802394, 2.1179683e-05, -3.5314584e-05, 1.8212895e-06, 7.693616e-07, -1.224184e-07, 0.0007326708, -2.5157635e-06, -3.4315726e-05, 2.483769e-06, 6.845847e-07, -1.3036272e-07, 0.00072561513, -2.5570285e-05, -3.2798627e-05, 3.0907177e-06, 5.90996e-07, -1.3604479e-07, 0.0007072656, -4.7635054e-05, -3.0800176e-05, 3.6338677e-06, 4.902957e-07, -1.3942868e-07, 0.0006781993, -6.838563e-05, -2.8363971e-05, 4.106167e-06, 3.8425554e-07, -1.4051592e-07, 0.0006391484, -8.7526496e-05, -2.5539486e-05, 4.501861e-06, 2.7468926e-07, -1.3934468e-07, 0.000590985, -0.00010479502, -2.2381117e-05, 4.8165534e-06, 1.6342224e-07, -1.359881e-07, 0.00053470343, -0.00011996482, -1.8947214e-05, 5.047241e-06, 5.2262546e-08, -1.3055244e-07, 0.00047140146, -0.00013284842, -1.529905e-05, 5.1923275e-06, -5.7027663e-08, -1.2317442e-07, 0.00040226066, -0.0001432993, -1.14997765e-05, 5.251616e-06, -1.6275894e-07, -1.1401841e-07, 0.00032852523, -0.00015121316, -7.613376e-06, 5.226276e-06, -2.6333964e-07, -1.0327305e-07, 0.00025148084, -0.0001565285, -3.7036243e-06, 5.1187903e-06, -3.5729894e-07, -9.1147704e-08, 0.00017243317, -0.00015922663, 1.6691529e-07, 4.932887e-06, -4.4330713e-07, -7.7868584e-08, 9.268676e-05, -0.0001593308, 3.937855e-06, 4.6734444e-06, -5.201934e-07, -6.3674754e-08, 1.3524288e-05, -0.00015690477, 7.5518883e-06, 4.34639e-06, -5.869605e-07, -4.8813988e-08, -6.3813175e-05, -0.00015205091, 1.0955622e-05, 3.9585775e-06, -6.4279635e-07, -3.3538637e-08, -0.00013814485, -0.0001449075, 1.4100328e-05, 3.5176565e-06, -6.870825e-07, -1.8101472e-08, -0.00020836745, -0.00013564568, 1.69426e-05, 3.0319297e-06, -7.19399e-07, -2.7516753e-09, -0.0002734707, -0.0001244659, 1.9444911e-05, 2.5102074e-06, -7.395264e-07, 1.22690595e-08, -0.0003325512, -0.000111594025, 2.1576061e-05, 1.9616527e-06, -7.4744423e-07, 2.6730177e-08, -0.0003848238, -9.72771e-05, 2.331152e-05, 1.3956285e-06, -7.433263e-07, 4.0415657e-08, -0.00042963136, -8.177891e-05, 2.4633646e-05, 8.2154384e-07, -7.275335e-07, 5.31271e-08, -0.00046645178, -6.537537e-05, 2.5531801e-05, 2.4870275e-07, -7.006031e-07, 6.468644e-08, -0.000494903, -4.8349815e-05, 2.6002335e-05, -3.138405e-07, -6.63236e-07, 7.4938285e-08, -0.0005147456, -3.0988376e-05, 2.6048481e-05, -8.5741925e-07, -6.162817e-07, 8.375184e-08, -0.0005258828, -1.3575309e-05, 2.5680129e-05, -1.3738822e-06, -5.607208e-07, 9.102237e-08, -0.0005283587, 3.6114407e-06, 2.49135e-05, -1.8557107e-06, -4.9764674e-07, 9.6672224e-08, -0.00052235374, 2.0304506e-05, 2.377073e-05, -2.2961217e-06, -4.2824496e-07, 1.006514e-07, -0.0005081787, 3.6251076e-05, 2.2279382e-05, -2.6891578e-06, -3.537724e-07, 1.02937676e-07, -0.0004862663, 5.121655e-05, 2.0471864e-05, -3.0297617e-06, -2.755354e-07, 1.0353629e-07, -0.00045716134, 6.49878e-05, 1.8384788e-05, -3.313833e-06, -1.9486785e-07, 1.0247913e-07, -0.00042150918, 7.737603e-05, 1.60583e-05, -3.5382716e-06, -1.131093e-07, 9.9823616e-08, -0.000380043, 8.821916e-05, 1.3535343e-05, -3.701e-06, -3.1583593e-08, 9.565116e-08, -0.00033356994, 9.738373e-05, 1.0860905e-05, -3.800972e-06, 4.842187e-08, 9.006524e-08, -0.00028295643, 0.00010476631, 8.081257e-06, -3.838164e-06, 1.2567561e-07, 8.318927e-08, -0.00022911289, 0.000110294386, 5.2431883e-06, -3.81355e-06, 1.9902028e-07, 7.5164095e-08, -0.00017297817, 0.00011392675, 2.3932444e-06, -3.7290602e-06, 2.673892e-07, 6.614533e-08, -0.00011550394, 0.00011565335, -4.2300243e-07, -3.5875275e-06, 3.2982112e-07, 5.6300575e-08, -5.76392e-05, 0.00011549469, -3.1616544e-06, -3.392621e-06, 3.8547276e-07, 4.580638e-08, -3.1529217e-07, 0.00011350073, -5.781143e-06, -3.1487652e-06, 4.336294e-07, 3.484528e-08, 5.5568486e-05, 0.00010974937, -8.242831e-06, -2.8610516e-06, 4.7371302e-07, 2.3602697e-08, 0.000109158354, 0.00010434448, -1.0511558e-05, -2.535142e-06, 5.052881e-07, 1.2263974e-08, 0.00015965852, 9.741363e-05, -1.2556102e-05, -2.1771634e-06, 5.2806485e-07, 1.011387e-09, 0.00020634232, 8.9105444e-05, -1.4349588e-05, -1.7935997e-06, 5.419006e-07, -9.978649e-09, 0.0002485621, 7.958674e-05, -1.5869802e-05, -1.3911796e-06, 5.4679793e-07, -2.053825e-08, 0.00028575756, 6.903941e-05, -1.7099426e-05, -9.767637e-07, 5.4290143e-07, -3.0510517e-08, 0.0003174623, 5.7657133e-05, -1.8026194e-05, -5.57232e-07, 5.3049166e-07, -3.975175e-08, 0.0003433092, 4.564202e-05, -1.8642962e-05, -1.3937465e-07, 5.099774e-07, -4.813342e-08, 0.00036303338, 3.320119e-05, -1.894769e-05, 2.7021417e-07, 4.818858e-07, -5.5543815e-08, 0.00037647423, 2.054335e-05, -1.8943347e-05, 6.65236e-07, 4.4685163e-07, -6.188942e-08, 0.00038357507, 7.875421e-06, -1.8637744e-05, 1.0397806e-06, 4.0560366e-07, -6.7095954e-08, 0.00038438165, -4.6006876e-06, -1.8043283e-05, 1.3884106e-06, 3.589515e-07, -7.110903e-08, 0.0003790387, -1.6691172e-05, -1.717665e-05, 1.7062358e-06, 3.0777036e-07, -7.389458e-08, 0.00036778528, -2.8213215e-05, -1.605844e-05, 1.9889774e-06, 2.5298564e-07, -7.5438884e-08, 0.00035094854, -3.8997616e-05, -1.4712734e-05, 2.2330203e-06, 1.955569e-07, -7.574824e-08, 0.00032893626, -4.8891143e-05, -1.3166626e-05, 2.435455e-06, 1.3646185e-07, -7.484843e-08, 0.00030222852, -5.7758567e-05, -1.1449722e-05, 2.594105e-06, 7.668032e-08, -7.278378e-08, 0.00027136807, -6.5484375e-05, -9.593601e-06, 2.7075446e-06, 1.7178682e-08, -6.9616014e-08, 0.00023695028, -7.19741e-05, -7.63127e-06, 2.7751014e-06, -4.110523e-08, -6.542285e-08, 0.00019961219, -7.715531e-05, -5.5965997e-06, 2.7968492e-06, -9.7276256e-08, -6.029636e-08, 0.00016002147, -8.097819e-05, -3.523763e-06, 2.7735878e-06, -1.5049508e-07, -5.4341136e-08, 0.000118865, -8.341581e-05, -1.4466889e-06, 2.7068122e-06, -1.9999023e-07, -4.767235e-08, 7.683738e-05, -8.446393e-05, 6.014751e-07, 2.5986722e-06, -2.4506852e-07, -4.041364e-08, 3.462978e-05, -8.4140534e-05, 2.5888683e-06, 2.4519204e-06, -2.8512426e-07, -3.269493e-08, -7.081018e-06, -8.2485e-05, 4.485392e-06, 2.2698553e-06, -3.1964666e-07, -2.4650234e-08, -4.764302e-05, -7.95569e-05, 6.2631434e-06, 2.0562536e-06, -3.482255e-07, -1.64154e-08, -8.6438784e-05, -7.5434575e-05, 7.896807e-06, 1.8152998e-06, -3.7055528e-07, -8.125928e-09, -0.00012289437, -7.0213435e-05, 9.363987e-06, 1.5515081e-06, -3.864373e-07, 8.51933e-11, -0.00015648743, -6.4003965e-05, 1.06455e-05, 1.2696436e-06, -3.957804e-07, 8.0895255e-09, -0.00018675414, -5.6929654e-05, 1.17255895e-05, 9.746391e-07, -3.9859947e-07, 1.576511e-08, -0.00021329525, -4.9124657e-05, 1.2592098e-05, 6.7151376e-07, -3.9501273e-07, 2.2998247e-08, -0.00023578072, -4.073142e-05, 1.3236568e-05, 3.652905e-07, -3.8523726e-07, 2.9685093e-08, -0.0002539533, -3.189819e-05, 1.3654284e-05, 6.091598e-08, -3.6958306e-07, 3.5733073e-08, -0.00026763082, -2.2776538e-05, 1.3844257e-05, -2.3681584e-07, -3.484458e-07, 4.1062062e-08, -0.00027670717, -1.3518837e-05, 1.3809143e-05, -5.2333627e-07, -3.2229843e-07, 4.5605354e-08, -0.00028115214, -4.275835e-06, 1.3555114e-05, -7.943688e-07, -2.9168174e-07, 4.9310387e-08, -0.00028100997, 4.8057086e-06, 1.3091668e-05, -1.04599e-06, -2.5719407e-07, 5.2139224e-08, -0.0002763968, 1.358526e-05, 1.24314e-05, -1.2746827e-06, -2.1948033e-07, 5.40688e-08, -0.00026749712, 2.1930588e-05, 1.1589721e-05, -1.4773825e-06, -1.792206e-07, 5.509091e-08, -0.000254559, 2.9719662e-05, 1.0584543e-05, -1.6515143e-06, -1.3711853e-07, 5.521197e-08, -0.0002378886, 3.684234e-05, 9.435933e-06, -1.7950216e-06, -9.388944e-08, 5.4452556e-08, -0.00021784393, 4.3201828e-05, 8.165739e-06, -1.9063863e-06, -5.0248765e-08, 5.2846726e-08, -0.00019482776, 4.871588e-05, 6.797201e-06, -1.9846393e-06, -6.900602e-09, 5.0441127e-08, -0.00016928017, 5.331775e-05, 5.354542e-06, -2.029362e-06, 3.5473143e-08, 4.729397e-08, -0.00014167058, 5.695687e-05, 3.862561e-06, -2.0406796e-06, 7.6223074e-08, 4.3473783e-08, -0.00011248953, 5.9599242e-05, 2.3462253e-06, -2.0192456e-06, 1.147418e-07, 3.905809e-08, -8.224043e-05, 6.1227576e-05, 8.30267e-07, -1.9662177e-06, 1.5047257e-07, 3.413195e-08, -5.143117e-05, 6.184115e-05, -6.6120367e-07, -1.8832275e-06, 1.8291682e-07, 2.878641e-08, -2.0565918e-05, 6.145541e-05, -2.1050662e-06, -1.772342e-06, 2.1164068e-07, 2.3116906e-08, 9.862763e-06, 6.0101294e-05, -3.4795332e-06, -1.6360209e-06, 2.3628027e-07, 1.7221655e-08, 3.9381503e-05, 5.7824407e-05, -4.7644635e-06, -1.4770666e-06, 2.565457e-07, 1.1200009e-08, 6.754316e-05, 5.4683886e-05, -5.9416407e-06, -1.298572e-06, 2.7222387e-07, 5.1508486e-09, 9.393329e-05, 5.0751136e-05, -6.995018e-06, -1.1038635e-06, 2.8317993e-07, -8.2897034e-10, 0.000118175914, 4.6108406e-05, -7.910915e-06, -8.9644243e-07, 2.8935747e-07, -6.64611e-09, 0.00013993857, 4.0847182e-05, -8.67818e-06, -6.799252e-07, 2.9077748e-07, -1.2212146e-08, 0.00015893648, 3.506652e-05, -9.288302e-06, -4.5798282e-07, 2.875361e-07, -1.7444851e-08};
	localparam real hb[0:1799] = {0.04146539, 0.00024480597, -0.00026783795, -2.248845e-06, 4.3801842e-06, 4.864713e-08, 0.041221026, 0.00073176116, -0.0002614101, -6.696438e-06, 4.290541e-06, 1.448581e-07, 0.040734954, 0.0012107815, -0.00024864986, -1.0994666e-05, 4.1132726e-06, 2.3784936e-07, 0.04001243, 0.0016766941, -0.0002297464, -1.5047003e-05, 3.8523635e-06, 3.2557224e-07, 0.039061278, 0.0021244998, -0.00020497982, -1.8761422e-05, 3.5136645e-06, 4.06118e-07, 0.037891746, 0.0025494383, -0.00017471658, -2.205205e-05, 3.1047541e-06, 4.7776365e-07, 0.036516394, 0.0029470513, -0.00013940375, -2.4840714e-05, 2.6347661e-06, 5.3901107e-07, 0.034949932, 0.0033132397, -9.9561985e-05, -2.7058317e-05, 2.1141852e-06, 5.8861855e-07, 0.03320901, 0.003644315, -5.5777306e-05, -2.8646065e-05, 1.5546185e-06, 6.256258e-07, 0.03131201, 0.003937048, -8.692036e-06, -2.9556486e-05, 9.685473e-07, 6.493704e-07, 0.029278811, 0.0041887052, 4.100521e-05, -2.9754228e-05, 3.690637e-07, 6.594982e-07, 0.027130522, 0.0043970835, 9.259013e-05, -2.9216664e-05, -2.3039931e-07, 6.559652e-07, 0.024889218, 0.0045605334, 0.00014531388, -2.7934244e-05, -8.163425e-07, 6.390335e-07, 0.02257766, 0.004677976, 0.00019841442, -2.5910616e-05, -1.3754711e-06, 6.092603e-07, 0.020218996, 0.0047489107, 0.00025112805, -2.3162525e-05, -1.8949582e-06, 5.6748127e-07, 0.01783649, 0.0047734166, 0.00030270085, -1.9719477e-05, -2.3626956e-06, 5.1478764e-07, 0.015453213, 0.0047521433, 0.00035239992, -1.5623187e-05, -2.7675267e-06, 4.5249982e-07, 0.013091778, 0.004686295, 0.00039952397, -1.0926819e-05, -3.0994586e-06, 3.8213585e-07, 0.010774061, 0.0045776074, 0.00044341368, -5.6940457e-06, -3.34985e-06, 3.053772e-07, 0.008520941, 0.004428317, 0.00048346096, 2.079197e-09, -3.5115697e-06, 2.2403161e-07, 0.0063520637, 0.004241123, 0.0005191175, 6.08038e-06, -3.579126e-06, 1.3999463e-07, 0.0042856177, 0.004019145, 0.0005499023, 1.2452956e-05, -3.548764e-06, 5.5209913e-08, 0.0023381365, 0.0037658734, 0.000575408, 1.902667e-05, -3.4185289e-06, -2.8370449e-08, 0.00052432675, 0.0034851169, 0.00059530616, 2.5704714e-05, -3.1882964e-06, -1.0882508e-07, -0.0011430768, 0.0031809455, 0.0006093511, 3.2388223e-05, -2.8597694e-06, -1.8430102e-07, -0.0026534274, 0.0028576308, 0.0006173824, 3.8977894e-05, -2.4364408e-06, -2.5304948e-07, -0.0039982516, 0.002519585, 0.0006193266, 4.5375622e-05, -1.9235256e-06, -3.1345897e-07, -0.0051713055, 0.0021712987, 0.00061519654, 5.1486055e-05, -1.3278617e-06, -3.640851e-07, -0.006168595, 0.0018172781, 0.0006050904, 5.721813e-05, -6.577848e-07, -4.036769e-07, -0.0069883717, 0.0014619845, 0.0005891891, 6.248652e-05, 7.702353e-08, -4.3119886e-07, -0.007631094, 0.001109774, 0.0005677523, 6.721291e-05, 8.65709e-07, -4.4584894e-07, -0.00809936, 0.0007648413, 0.00054111326, 7.132724e-05, 1.6964362e-06, -4.4707144e-07, -0.008397813, 0.00043116606, 0.00050967326, 7.476873e-05, 2.5565953e-06, -4.345657e-07, -0.008533023, 0.000112463655, 0.00047389444, 7.748676e-05, 3.43302e-06, -4.0828954e-07, -0.008513342, -0.00018785929, 0.00043429201, 7.9441576e-05, 4.3122127e-06, -3.684583e-07, -0.008348739, -0.00046674386, 0.00039142597, 8.0604856e-05, 5.180572e-06, -3.1553893e-07, -0.00805062, -0.00072151225, 0.00034589216, 8.096e-05, 6.0246216e-06, -2.5023982e-07, -0.007631627, -0.0009498948, 0.000298313, 8.05023e-05, 6.831232e-06, -1.7349653e-07, -0.007105432, -0.0011500503, 0.00024932786, 7.923891e-05, 7.5878356e-06, -8.645332e-08, -0.0064865164, -0.0013205807, 0.00019958348, 7.71886e-05, 8.282629e-06, 9.558333e-09, -0.0057899496, -0.0014605374, 0.00014972452, 7.4381336e-05, 8.904762e-06, 1.1304449e-07, -0.00503116, -0.001569423, 0.00010038412, 7.085774e-05, 9.444505e-06, 2.2237596e-07, -0.004225716, -0.0016471844, 5.217493e-05, 6.6668326e-05, 9.893401e-06, 3.3581745e-07, -0.0033891022, -0.0016942013, 5.6806734e-06, 6.187262e-05, 1.0244392e-05, 4.5155824e-07, -0.0025365087, -0.0017112679, -3.8551792e-05, 5.6538138e-05, 1.0491919e-05, 5.6774377e-07, -0.0016826305, -0.0016995692, -8.001964e-05, 5.07393e-05, 1.0632002e-05, 6.825074e-07, -0.0008414778, -0.0016606523, -0.00011827045, 4.4556207e-05, 1.06622865e-05, 7.9400235e-07, -2.6203514e-05, -0.0015963936, -0.0001529077, 3.807334e-05, 1.0582069e-05, 9.0043227e-07, 0.00075105205, -0.0015089608, -0.00018359527, 3.1378277e-05, 1.0392294e-05, 1.0000812e-06, 0.0014792971, -0.0014007733, -0.00021006101, 2.4560304e-05, 1.009552e-05, 1.0913416e-06, 0.002148803, -0.0012744586, -0.00023209922, 1.7709088e-05, 9.695872e-06, 1.1727395e-06, 0.0027511988, -0.0011328079, -0.00024957207, 1.0913319e-05, 9.1989505e-06, 1.2429585e-06, 0.0032795395, -0.0009787299, -0.00026241003, 4.2594206e-06, 8.61174e-06, 1.3008598e-06, 0.0037283541, -0.0008152043, -0.00027061123, -2.169698e-06, 7.942478e-06, 1.3454986e-06, 0.00409367, -0.0006452354, -0.00027423972, -8.295808e-06, 7.2005223e-06, 1.3761386e-06, 0.0043730135, -0.0004718075, -0.00027342307, -1.4046433e-05, 6.396189e-06, 1.3922617e-06, 0.004565388, -0.00029784048, -0.00026834864, -1.935582e-05, 5.5405853e-06, 1.393574e-06, 0.0046712337, -0.00012614891, -0.00025925948, -2.4165789e-05, 4.645431e-06, 1.3800093e-06, 0.004692362, 4.059674e-05, -0.0002464492, -2.8426433e-05, 3.7228735e-06, 1.3517264e-06, 0.004631878, 0.00019990538, -0.00023025631, -3.2096712e-05, 2.785297e-06, 1.3091061e-06, 0.004494078, 0.0003494969, -0.00021105794, -3.514487e-05, 1.8451333e-06, 1.2527415e-06, 0.0042843423, 0.0004873296, -0.0001892633, -3.7548714e-05, 9.1467405e-07, 1.1834273e-06, 0.004009006, 0.0006116232, -0.00016530664, -3.929575e-05, 5.888459e-09, 1.1021446e-06, 0.003675227, 0.0007208773, -0.00013964009, -4.038316e-05, -8.697514e-07, 1.0100435e-06, 0.0032908383, 0.0008138848, -0.00011272643, -4.0817617e-05, -1.701434e-06, 9.08424e-07, 0.0028642027, 0.0008897404, -8.5031825e-05, -4.0615e-05, -2.4791593e-06, 7.9871296e-07, 0.0024040581, 0.00094784505, -5.701874e-05, -3.9799936e-05, -3.1938737e-06, 6.8244145e-07, 0.0019193669, 0.0009879041, -2.9139079e-05, -3.8405236e-05, -3.837589e-06, 5.6121934e-07, 0.0014191625, 0.0010099224, -1.8276651e-06, -3.647122e-05, -4.4034823e-06, 4.367096e-07, 0.0009124039, 0.0010141934, 2.450384e-05, -3.4044948e-05, -4.885976e-06, 3.1060247e-07, 0.00040783366, 0.0010012859, 4.9472517e-05, -3.1179337e-05, -5.2807973e-06, 1.845891e-07, -8.6154956e-05, 0.00097202475, 7.272916e-05, -2.793225e-05, -5.585017e-06, 6.033577e-08, -0.000561641, 0.0009274706, 9.396263e-05, -2.4365498e-05, -5.797066e-06, -6.0540856e-08, -0.0010112876, 0.0008688947, 0.000112903464, -2.0543823e-05, -5.916733e-06, -1.7649754e-07, -0.0014284403, 0.0007977517, 0.00012932679, -1.6533855e-05, -5.9451363e-06, -2.8608656e-07, -0.0018072124, 0.00071565114, 0.00014305445, -1.240306e-05, -5.884684e-06, -3.8797606e-07, -0.0021425537, 0.0006243265, 0.00015395635, -8.218712e-06, -5.7390066e-06, -4.809681e-07, -0.0024303054, 0.00052560354, 0.00016195106, -4.046875e-06, -5.5128776e-06, -5.640142e-07, -0.0026672382, 0.00042136834, 0.00016700556, 4.855194e-08, -5.212119e-06, -6.36229e-07, -0.002851074, 0.0003135352, 0.00016913444, 4.006748e-06, -4.8434886e-06, -6.9689986e-07, -0.0029804923, 0.00020401487, 0.00016839804, 7.770807e-06, -4.4145577e-06, -7.454949e-07, -0.0030551208, 9.468427e-05, 0.00016490035, 1.1288498e-05, -3.9335814e-06, -7.816673e-07, -0.0030755112, -1.2642788e-05, 0.00015878597, 1.451293e-05, -3.4093562e-06, -8.05257e-07, -0.0030431, -0.000116242794, 0.00015023665, 1.7403117e-05, -2.8510776e-06, -8.162893e-07, -0.0029601583, -0.00021450751, 0.00013946736, 1.9924453e-05, -2.2681913e-06, -8.1497086e-07, -0.0028297275, -0.0003059664, 0.00012672189, 2.2049056e-05, -1.6702459e-06, -8.0168275e-07, -0.002655546, -0.0003893061, 0.0001122682, 2.3756009e-05, -1.066746e-06, -7.769712e-07, -0.0024419657, -0.00046338706, 9.639343e-05, 2.5031492e-05, -4.6701115e-07, -7.415358e-07, -0.002193862, -0.0005272565, 7.939882e-05, 2.58688e-05, 1.1996097e-07, -6.9621575e-07, -0.0019165382, -0.00058015855, 6.159456e-05, 2.6268237e-05, 6.856217e-07, -6.4197405e-07, -0.0016156246, -0.00062154036, 4.3294538e-05, 2.6236929e-05, 1.2219896e-06, -5.798804e-07, -0.0012969768, -0.00065105513, 2.4811325e-05, 2.578851e-05, 1.7217562e-06, -5.1109276e-07, -0.00096657197, -0.0006685619, 6.4511933e-06, 2.4942734e-05, 2.1783806e-06, -4.368377e-07, -0.0006304072, -0.0006741216, -1.1490546e-05, 2.3725e-05, 2.5861673e-06, -3.5839042e-07, -0.00029439994, -0.0006679901, -2.8733944e-05, 2.2165796e-05, 2.9403316e-06, -2.770545e-07, 3.570702e-05, -0.00065060885, -4.5018438e-05, 2.030007e-05, 3.2370483e-06, -1.9414136e-07, 0.0003544354, -0.00062259194, -6.0106442e-05, 1.8166582e-05, 3.4734844e-06, -1.10950424e-07, 0.0006566542, -0.00058471126, -7.378651e-05, 1.580717e-05, 3.6478157e-06, -2.8749648e-08, 0.0009376542, -0.0005378797, -8.587597e-05, 1.32660225e-05, 3.759228e-06, 5.124282e-08, 0.001193214, -0.0004831321, -9.6223e-05, 1.0588912e-05, 3.8079017e-06, 1.2787592e-07, 0.0014196559, -0.00042160501, -0.00010470825, 7.822441e-06, 3.794983e-06, 2.0008146e-07, 0.0016138916, -0.0003545153, -0.000111245805, 5.0132785e-06, 3.7225384e-06, 2.668882e-07, 0.0017734565, -0.0002831382, -0.000115783645, 2.2074303e-06, 3.5934993e-06, 3.2743432e-07, 0.0018965335, -0.00020878478, -0.00011830353, -5.504701e-07, 3.411592e-06, 3.8097758e-07, 0.001981966, -0.00013277972, -0.000118820346, -3.2178243e-06, 3.1812583e-06, 4.269036e-07, 0.0020292576, -5.6439232e-05, -0.000117380994, -5.7546863e-06, 2.907567e-06, 4.6473204e-07, 0.002038564, 1.895013e-05, -0.00011406272, -8.124317e-06, 2.5961187e-06, 4.941203e-07, 0.0020106724, 9.2151655e-05, -0.00010897106, -1.0293679e-05, 2.2529423e-06, 5.148652e-07, 0.0019469721, 0.0001619973, -0.00010223735, -1.2233855e-05, 1.8843914e-06, 5.269025e-07, 0.0018494154, 0.00022740495, -9.401595e-05, -1.3920389e-05, 1.4970343e-06, 5.3030413e-07, 0.001720471, 0.00028739372, -8.448112e-05, -1.5333557e-05, 1.097547e-06, 5.252735e-07, 0.0015630699, 0.0003410973, -7.382368e-05, -1.6458544e-05, 6.926051e-07, 5.121386e-07, 0.0013805453, 0.00038777513, -6.22475e-05, -1.7285545e-05, 2.887793e-07, 4.9134405e-07, 0.0011765675, 0.00042682106, -4.9965845e-05, -1.7809787e-05, -1.0756439e-07, 4.6344078e-07, 0.0009550746, 0.0004577699, -3.719775e-05, -1.803146e-05, -4.90359e-07, 4.2907462e-07, 0.00072020135, 0.00048030124, -2.4164285e-05, -1.7955588e-05, -8.539238e-07, 3.8897377e-07, 0.00047620616, 0.0004942409, -1.10849605e-05, -1.7591809e-05, -1.1930427e-06, 3.4393543e-07, 0.000227398, 0.0004995602, 1.8257559e-06, -1.6954098e-05, -1.503034e-06, 2.9481123e-07, -2.1935415e-05, 0.0004963725, 1.4361768e-05, -1.6060432e-05, -1.7798089e-06, 2.4249272e-07, -0.0002675976, 0.00048492796, 2.6328446e-05, -1.4932386e-05, -2.0199202e-06, 1.8789628e-07, -0.0005055498, 0.00046560587, 3.7545466e-05, -1.35947e-05, -2.2205988e-06, 1.3194817e-07, -0.0007319731, 0.00043890523, 4.7849324e-05, -1.2074796e-05, -2.379779e-06, 7.556981e-08, -0.000943326, 0.0004054338, 5.7095556e-05, -1.0402267e-05, -2.496112e-06, 1.966345e-08, -0.0011363953, 0.00036589528, 6.516055e-05, -8.608349e-06, -2.5689671e-06, -3.490142e-08, -0.0013083407, 0.00032107567, 7.194299e-05, -6.7253745e-06, -2.5984232e-06, -8.7300805e-08, -0.0014567326, 0.0002718284, 7.736494e-05, -4.7862313e-06, -2.585247e-06, -1.3676791e-07, -0.0015795819, 0.00021905889, 8.1372455e-05, -2.823819e-06, -2.5308632e-06, -1.8260363e-07, -0.0016753613, 0.00016370844, 8.393588e-05, -8.705237e-07, -2.4373128e-06, -2.2418568e-07, -0.0017430203, 0.00010673826, 8.504967e-05, 1.0422855e-06, -2.3072055e-06, -2.6097635e-07, -0.0017819905, 4.9113318e-05, 8.473187e-05, 2.884732e-06, -2.1436617e-06, -2.9252863e-07, -0.0017921835, -8.213343e-06, 8.302324e-05, 4.62887e-06, -1.9502497e-06, -3.184908e-07, -0.0017739814, -6.431576e-05, 7.998597e-05, 6.249081e-06, -1.7309167e-06, -3.386095e-07, -0.0017282194, -0.00011830935, 7.5702206e-05, 7.7224195e-06, -1.4899155e-06, -3.527309e-07, -0.0016561622, -0.00016936421, 7.027217e-05, 9.028916e-06, -1.2317291e-06, -3.6080053e-07, -0.0015594726, -0.00021671722, 6.381213e-05, 1.0151813e-05, -9.609931e-07, -3.6286144e-07, -0.0014401767, -0.00025968274, 5.6452052e-05, 1.1077749e-05, -6.824175e-07, -3.5905097e-07, -0.0013006215, -0.00029766184, 4.8333266e-05, 1.1796891e-05, -4.0070975e-07, -3.4959587e-07, -0.0011434306, -0.00033014987, 3.9605828e-05, 1.230299e-05, -1.2049978e-07, -3.3480643e-07, -0.00097145484, -0.0003567423, 3.0425923e-05, 1.2593396e-05, 1.537317e-07, -3.150693e-07, -0.00078772154, -0.00037713893, 2.0953192e-05, 1.2668999e-05, 4.1772083e-07, -2.9083918e-07, -0.0005953814, -0.0003911462, 1.134808e-05, 1.2534132e-05, 6.6748277e-07, -2.6263004e-07, -0.00039765524, -0.00039867766, 1.7692399e-06, 1.2196404e-05, 8.99368e-07, -2.3100505e-07, -0.00019778035, -0.00039975307, -7.628977e-06, 1.1666498e-05, 1.1101118e-06, -1.965666e-07, 1.0417496e-06, -0.00039449532, -1.669889e-05, 1.0957918e-05, 1.296876e-06, -1.599455e-07, 0.00019569589, -0.0003831261, -2.5301697e-05, 1.0086704e-05, 1.4572834e-06, -1.2179028e-07, 0.00038320126, -0.00036596006, -3.3309487e-05, 9.071102e-06, 1.5894433e-06, -8.275637e-08, 0.0005607561, -0.00034339743, -4.0607014e-05, 7.931223e-06, 1.6919691e-06, -4.349549e-08, 0.00072577846, -0.00031591573, -4.709325e-05, 6.6886664e-06, 1.7639875e-06, -4.645376e-09, 0.0008759425, -0.0002840602, -5.2682648e-05, 5.3661397e-06, 1.8051384e-06, 3.3179994e-08, 0.0010092098, -0.0002484334, -5.7306126e-05, 3.987063e-06, 1.8155679e-06, 6.939956e-08, 0.0011238554, -0.00020968445, -6.091179e-05, 2.5751765e-06, 1.7959125e-06, 1.0347359e-07, 0.0012184877, -0.00016849731, -6.346532e-05, 1.1541526e-06, 1.7472757e-06, 1.3491113e-07, 0.0012920641, -0.00012557908, -6.4950116e-05, -2.5278408e-07, 1.6711991e-06, 1.6327662e-07, 0.0013438981, -8.164823e-05, -6.5367116e-05, -1.623217e-06, 1.5696256e-06, 1.8819536e-07, 0.0013736633, -3.742277e-05, -6.473434e-05, -2.9358766e-06, 1.4448581e-06, 2.0935782e-07, 0.0013813896, 6.3911475e-06, -6.308622e-05, -4.170953e-06, 1.2995133e-06, 2.26523e-07, 0.0013674548, 4.9110262e-05, -6.047262e-05, -5.310377e-06, 1.136472e-06, 2.3952038e-07, 0.0013325703, 9.008453e-05, -5.695766e-05, -6.3380653e-06, 9.588255e-07, 2.4825076e-07, 0.0012777626, 0.00012870673, -5.261836e-05, -7.24013e-06, 7.6982104e-07, 2.5268616e-07, 0.0012043486, 0.00016442109, -4.7543097e-05, -8.005044e-06, 5.7280613e-07, 2.528682e-07, 0.0011139092, 0.00019673095, -4.182989e-05, -8.623769e-06, 3.7117152e-07, 2.4890576e-07, 0.0010082573, 0.00022520528, -3.558463e-05, -9.089839e-06, 1.6829631e-07, 2.4097142e-07, 0.00088940363, 0.00024948397, -2.8919168e-05, -9.399396e-06, -3.250605e-08, 2.2929709e-07, 0.00075952057, 0.00026928185, -2.1949405e-05, -9.5511905e-06, -2.2803921e-07, 2.1416871e-07, 0.0006209036, 0.00028439148, -1.4793331e-05, -9.546537e-06, -4.1527218e-07, 1.9592031e-07, 0.00047593226, 0.00029468464, -7.569097e-06, -9.389224e-06, -5.9138364e-07, 1.7492742e-07, 0.0003270303, 0.00030011236, -3.9312047e-07, -9.0854e-06, -7.5380206e-07, 1.5160002e-07, 0.00017662637, 0.0003007039, 6.621728e-06, -8.643411e-06, -9.002402e-07, 1.2637503e-07, 2.7115331e-05, 0.00029656442, 1.3367841e-05, -8.073614e-06, -1.0287251e-06, 9.970865e-08, -0.000119178745, 0.00028787146, 1.9744464e-05, -7.3881624e-06, -1.1376214e-06, 7.206857e-08, -0.00026003775, 0.0002748704, 2.565913e-05, -6.6007674e-06, -1.2256492e-06, 4.392621e-08, -0.0003933821, 0.00025786896, 3.1028943e-05, -5.7264383e-06, -1.2918955e-06, 1.5749015e-08, -0.00051730033, 0.0002372308, 3.5781653e-05, -4.7812127e-06, -1.3358201e-06, -1.2006875e-08, -0.0006300753, 0.00021336837, 3.9856568e-05, -3.781874e-06, -1.3572542e-06, -3.890365e-08, -0.0007302067, 0.0001867353, 4.320522e-05, -2.7456647e-06, -1.3563944e-06, -6.452839e-08, -0.00081642973, 0.00015781808, 4.5791854e-05, -1.6899994e-06, -1.3337901e-06, -8.849904e-08, -0.00088772917, 0.00012712766, 4.759369e-05, -6.3218243e-07, -1.2903263e-06, -1.10469735e-07, -0.0009433496, 9.51907e-05, 4.8600963e-05, 4.108655e-07, -1.2272005e-06, -1.3013542e-07, -0.0009828011, 6.254085e-05, 4.881676e-05, 1.4228688e-06, -1.1458965e-06, -1.4723571e-07, -0.0010058604, 2.9710145e-05, 4.8256672e-05, 2.3884404e-06, -1.0481527e-06, -1.6155796e-07, -0.0010125681, -2.7794342e-06, 4.6948237e-05, 3.2933067e-06, -9.359288e-07, -1.7293941e-07, -0.001003222, -3.4423952e-05, 4.49302e-05, 4.124507e-06, -8.1136835e-07, -1.8126859e-07, -0.000978365, -6.474508e-05, 4.225164e-05, 4.870569e-06, -6.767601e-07, -1.8648575e-07, -0.00093877193, -9.3297065e-05, 3.8970928e-05, 5.521654e-06, -5.344981e-07, -1.885826e-07, -0.00088543084, -0.000119672986, 3.5154586e-05, 6.0696775e-06, -3.870403e-07, -1.8760112e-07, -0.0008195223, -0.00014351026, 3.0876014e-05, 6.508391e-06, -2.3686813e-07, -1.8363157e-07, -0.0007423962, -0.0001644953, 2.6214162e-05, 6.833439e-06, -8.644602e-08, -1.7680995e-07, -0.00065554614, -0.00018236731, 2.1252148e-05, 7.0423816e-06, 6.181753e-08, -1.6731461e-07, -0.00056058227, -0.00019692112, 1.6075826e-05, 7.134687e-06, 2.0560704e-07, -1.5536234e-07, -0.000459203, -0.00020800902, 1.0772361e-05, 7.111694e-06, 3.427347e-07, -1.4120398e-07, -0.0003531661, -0.00021554178, 5.4288053e-06, 6.976542e-06, 4.7117229e-07, -1.2511956e-07, -0.00024425922, -0.00021948859, 1.3072744e-07, 6.734081e-06, 5.890795e-07, -1.0741304e-07, -0.00013427105, -0.00021987609, -5.0391163e-06, 6.39075e-06, 6.948289e-07, -8.840692e-08, -2.4962921e-05, -0.0002167866, -1.0002027e-05, 5.954436e-06, 7.870264e-07, -6.843662e-08, 8.195832e-05, -0.00021035537, -1.46845105e-05, 5.434313e-06, 8.645281e-07, -4.7844743e-08, 0.00018486603, -0.0002007672, -1.901932e-05, 4.8406664e-06, 9.264522e-07, -2.6975489e-08, 0.00028223748, -0.00018825223, -2.2946373e-05, 4.184698e-06, 9.721866e-07, -6.1690666e-09, 0.0003726754, -0.00017308127, -2.641352e-05, 3.4783302e-06, 1.0013924e-06, 1.4243616e-08, 0.00045492692, -0.00015556037, -2.9377186e-05, 2.7339945e-06, 1.0140021e-06, 3.394602e-08, 0.00052789995, -0.00013602525, -3.1802854e-05, 1.964424e-06, 1.0102143e-06, 5.2640676e-08, 0.00059067627, -0.00011483514, -3.3665376e-05, 1.1824418e-06, 9.904842e-07, 7.005346e-08, 0.00064252195, -9.236654e-05, -3.4949164e-05, 4.0075614e-07, 9.555097e-07, 8.5937394e-08, 0.00068289426, -6.900684e-05, -3.564818e-05, -3.6824008e-07, 9.0621444e-07, 1.0007594e-07, 0.0007114456, -4.5147888e-05, -3.5765814e-05, -1.112658e-06, 8.4372783e-07, 1.1228567e-07, 0.00072802394, -2.1179683e-05, -3.5314584e-05, -1.8212895e-06, 7.693616e-07, 1.224184e-07, 0.0007326708, 2.5157635e-06, -3.4315726e-05, -2.483769e-06, 6.845847e-07, 1.3036272e-07, 0.00072561513, 2.5570285e-05, -3.2798627e-05, -3.0907177e-06, 5.90996e-07, 1.3604479e-07, 0.0007072656, 4.7635054e-05, -3.0800176e-05, -3.6338677e-06, 4.902957e-07, 1.3942868e-07, 0.0006781993, 6.838563e-05, -2.8363971e-05, -4.106167e-06, 3.8425554e-07, 1.4051592e-07, 0.0006391484, 8.7526496e-05, -2.5539486e-05, -4.501861e-06, 2.7468926e-07, 1.3934468e-07, 0.000590985, 0.00010479502, -2.2381117e-05, -4.8165534e-06, 1.6342224e-07, 1.359881e-07, 0.00053470343, 0.00011996482, -1.8947214e-05, -5.047241e-06, 5.2262546e-08, 1.3055244e-07, 0.00047140146, 0.00013284842, -1.529905e-05, -5.1923275e-06, -5.7027663e-08, 1.2317442e-07, 0.00040226066, 0.0001432993, -1.14997765e-05, -5.251616e-06, -1.6275894e-07, 1.1401841e-07, 0.00032852523, 0.00015121316, -7.613376e-06, -5.226276e-06, -2.6333964e-07, 1.0327305e-07, 0.00025148084, 0.0001565285, -3.7036243e-06, -5.1187903e-06, -3.5729894e-07, 9.1147704e-08, 0.00017243317, 0.00015922663, 1.6691529e-07, -4.932887e-06, -4.4330713e-07, 7.7868584e-08, 9.268676e-05, 0.0001593308, 3.937855e-06, -4.6734444e-06, -5.201934e-07, 6.3674754e-08, 1.3524288e-05, 0.00015690477, 7.5518883e-06, -4.34639e-06, -5.869605e-07, 4.8813988e-08, -6.3813175e-05, 0.00015205091, 1.0955622e-05, -3.9585775e-06, -6.4279635e-07, 3.3538637e-08, -0.00013814485, 0.0001449075, 1.4100328e-05, -3.5176565e-06, -6.870825e-07, 1.8101472e-08, -0.00020836745, 0.00013564568, 1.69426e-05, -3.0319297e-06, -7.19399e-07, 2.7516753e-09, -0.0002734707, 0.0001244659, 1.9444911e-05, -2.5102074e-06, -7.395264e-07, -1.22690595e-08, -0.0003325512, 0.000111594025, 2.1576061e-05, -1.9616527e-06, -7.4744423e-07, -2.6730177e-08, -0.0003848238, 9.72771e-05, 2.331152e-05, -1.3956285e-06, -7.433263e-07, -4.0415657e-08, -0.00042963136, 8.177891e-05, 2.4633646e-05, -8.2154384e-07, -7.275335e-07, -5.31271e-08, -0.00046645178, 6.537537e-05, 2.5531801e-05, -2.4870275e-07, -7.006031e-07, -6.468644e-08, -0.000494903, 4.8349815e-05, 2.6002335e-05, 3.138405e-07, -6.63236e-07, -7.4938285e-08, -0.0005147456, 3.0988376e-05, 2.6048481e-05, 8.5741925e-07, -6.162817e-07, -8.375184e-08, -0.0005258828, 1.3575309e-05, 2.5680129e-05, 1.3738822e-06, -5.607208e-07, -9.102237e-08, -0.0005283587, -3.6114407e-06, 2.49135e-05, 1.8557107e-06, -4.9764674e-07, -9.6672224e-08, -0.00052235374, -2.0304506e-05, 2.377073e-05, 2.2961217e-06, -4.2824496e-07, -1.006514e-07, -0.0005081787, -3.6251076e-05, 2.2279382e-05, 2.6891578e-06, -3.537724e-07, -1.02937676e-07, -0.0004862663, -5.121655e-05, 2.0471864e-05, 3.0297617e-06, -2.755354e-07, -1.0353629e-07, -0.00045716134, -6.49878e-05, 1.8384788e-05, 3.313833e-06, -1.9486785e-07, -1.0247913e-07, -0.00042150918, -7.737603e-05, 1.60583e-05, 3.5382716e-06, -1.131093e-07, -9.9823616e-08, -0.000380043, -8.821916e-05, 1.3535343e-05, 3.701e-06, -3.1583593e-08, -9.565116e-08, -0.00033356994, -9.738373e-05, 1.0860905e-05, 3.800972e-06, 4.842187e-08, -9.006524e-08, -0.00028295643, -0.00010476631, 8.081257e-06, 3.838164e-06, 1.2567561e-07, -8.318927e-08, -0.00022911289, -0.000110294386, 5.2431883e-06, 3.81355e-06, 1.9902028e-07, -7.5164095e-08, -0.00017297817, -0.00011392675, 2.3932444e-06, 3.7290602e-06, 2.673892e-07, -6.614533e-08, -0.00011550394, -0.00011565335, -4.2300243e-07, 3.5875275e-06, 3.2982112e-07, -5.6300575e-08, -5.76392e-05, -0.00011549469, -3.1616544e-06, 3.392621e-06, 3.8547276e-07, -4.580638e-08, -3.1529217e-07, -0.00011350073, -5.781143e-06, 3.1487652e-06, 4.336294e-07, -3.484528e-08, 5.5568486e-05, -0.00010974937, -8.242831e-06, 2.8610516e-06, 4.7371302e-07, -2.3602697e-08, 0.000109158354, -0.00010434448, -1.0511558e-05, 2.535142e-06, 5.052881e-07, -1.2263974e-08, 0.00015965852, -9.741363e-05, -1.2556102e-05, 2.1771634e-06, 5.2806485e-07, -1.011387e-09, 0.00020634232, -8.9105444e-05, -1.4349588e-05, 1.7935997e-06, 5.419006e-07, 9.978649e-09, 0.0002485621, -7.958674e-05, -1.5869802e-05, 1.3911796e-06, 5.4679793e-07, 2.053825e-08, 0.00028575756, -6.903941e-05, -1.7099426e-05, 9.767637e-07, 5.4290143e-07, 3.0510517e-08, 0.0003174623, -5.7657133e-05, -1.8026194e-05, 5.57232e-07, 5.3049166e-07, 3.975175e-08, 0.0003433092, -4.564202e-05, -1.8642962e-05, 1.3937465e-07, 5.099774e-07, 4.813342e-08, 0.00036303338, -3.320119e-05, -1.894769e-05, -2.7021417e-07, 4.818858e-07, 5.5543815e-08, 0.00037647423, -2.054335e-05, -1.8943347e-05, -6.65236e-07, 4.4685163e-07, 6.188942e-08, 0.00038357507, -7.875421e-06, -1.8637744e-05, -1.0397806e-06, 4.0560366e-07, 6.7095954e-08, 0.00038438165, 4.6006876e-06, -1.8043283e-05, -1.3884106e-06, 3.589515e-07, 7.110903e-08, 0.0003790387, 1.6691172e-05, -1.717665e-05, -1.7062358e-06, 3.0777036e-07, 7.389458e-08, 0.00036778528, 2.8213215e-05, -1.605844e-05, -1.9889774e-06, 2.5298564e-07, 7.5438884e-08, 0.00035094854, 3.8997616e-05, -1.4712734e-05, -2.2330203e-06, 1.955569e-07, 7.574824e-08, 0.00032893626, 4.8891143e-05, -1.3166626e-05, -2.435455e-06, 1.3646185e-07, 7.484843e-08, 0.00030222852, 5.7758567e-05, -1.1449722e-05, -2.594105e-06, 7.668032e-08, 7.278378e-08, 0.00027136807, 6.5484375e-05, -9.593601e-06, -2.7075446e-06, 1.7178682e-08, 6.9616014e-08, 0.00023695028, 7.19741e-05, -7.63127e-06, -2.7751014e-06, -4.110523e-08, 6.542285e-08, 0.00019961219, 7.715531e-05, -5.5965997e-06, -2.7968492e-06, -9.7276256e-08, 6.029636e-08, 0.00016002147, 8.097819e-05, -3.523763e-06, -2.7735878e-06, -1.5049508e-07, 5.4341136e-08, 0.000118865, 8.341581e-05, -1.4466889e-06, -2.7068122e-06, -1.9999023e-07, 4.767235e-08, 7.683738e-05, 8.446393e-05, 6.014751e-07, -2.5986722e-06, -2.4506852e-07, 4.041364e-08, 3.462978e-05, 8.4140534e-05, 2.5888683e-06, -2.4519204e-06, -2.8512426e-07, 3.269493e-08, -7.081018e-06, 8.2485e-05, 4.485392e-06, -2.2698553e-06, -3.1964666e-07, 2.4650234e-08, -4.764302e-05, 7.95569e-05, 6.2631434e-06, -2.0562536e-06, -3.482255e-07, 1.64154e-08, -8.6438784e-05, 7.5434575e-05, 7.896807e-06, -1.8152998e-06, -3.7055528e-07, 8.125928e-09, -0.00012289437, 7.0213435e-05, 9.363987e-06, -1.5515081e-06, -3.864373e-07, -8.51933e-11, -0.00015648743, 6.4003965e-05, 1.06455e-05, -1.2696436e-06, -3.957804e-07, -8.0895255e-09, -0.00018675414, 5.6929654e-05, 1.17255895e-05, -9.746391e-07, -3.9859947e-07, -1.576511e-08, -0.00021329525, 4.9124657e-05, 1.2592098e-05, -6.7151376e-07, -3.9501273e-07, -2.2998247e-08, -0.00023578072, 4.073142e-05, 1.3236568e-05, -3.652905e-07, -3.8523726e-07, -2.9685093e-08, -0.0002539533, 3.189819e-05, 1.3654284e-05, -6.091598e-08, -3.6958306e-07, -3.5733073e-08, -0.00026763082, 2.2776538e-05, 1.3844257e-05, 2.3681584e-07, -3.484458e-07, -4.1062062e-08, -0.00027670717, 1.3518837e-05, 1.3809143e-05, 5.2333627e-07, -3.2229843e-07, -4.5605354e-08, -0.00028115214, 4.275835e-06, 1.3555114e-05, 7.943688e-07, -2.9168174e-07, -4.9310387e-08, -0.00028100997, -4.8057086e-06, 1.3091668e-05, 1.04599e-06, -2.5719407e-07, -5.2139224e-08, -0.0002763968, -1.358526e-05, 1.24314e-05, 1.2746827e-06, -2.1948033e-07, -5.40688e-08, -0.00026749712, -2.1930588e-05, 1.1589721e-05, 1.4773825e-06, -1.792206e-07, -5.509091e-08, -0.000254559, -2.9719662e-05, 1.0584543e-05, 1.6515143e-06, -1.3711853e-07, -5.521197e-08, -0.0002378886, -3.684234e-05, 9.435933e-06, 1.7950216e-06, -9.388944e-08, -5.4452556e-08, -0.00021784393, -4.3201828e-05, 8.165739e-06, 1.9063863e-06, -5.0248765e-08, -5.2846726e-08, -0.00019482776, -4.871588e-05, 6.797201e-06, 1.9846393e-06, -6.900602e-09, -5.0441127e-08, -0.00016928017, -5.331775e-05, 5.354542e-06, 2.029362e-06, 3.5473143e-08, -4.729397e-08, -0.00014167058, -5.695687e-05, 3.862561e-06, 2.0406796e-06, 7.6223074e-08, -4.3473783e-08, -0.00011248953, -5.9599242e-05, 2.3462253e-06, 2.0192456e-06, 1.147418e-07, -3.905809e-08, -8.224043e-05, -6.1227576e-05, 8.30267e-07, 1.9662177e-06, 1.5047257e-07, -3.413195e-08, -5.143117e-05, -6.184115e-05, -6.6120367e-07, 1.8832275e-06, 1.8291682e-07, -2.878641e-08, -2.0565918e-05, -6.145541e-05, -2.1050662e-06, 1.772342e-06, 2.1164068e-07, -2.3116906e-08, 9.862763e-06, -6.0101294e-05, -3.4795332e-06, 1.6360209e-06, 2.3628027e-07, -1.7221655e-08, 3.9381503e-05, -5.7824407e-05, -4.7644635e-06, 1.4770666e-06, 2.565457e-07, -1.1200009e-08, 6.754316e-05, -5.4683886e-05, -5.9416407e-06, 1.298572e-06, 2.7222387e-07, -5.1508486e-09, 9.393329e-05, -5.0751136e-05, -6.995018e-06, 1.1038635e-06, 2.8317993e-07, 8.2897034e-10, 0.000118175914, -4.6108406e-05, -7.910915e-06, 8.9644243e-07, 2.8935747e-07, 6.64611e-09, 0.00013993857, -4.0847182e-05, -8.67818e-06, 6.799252e-07, 2.9077748e-07, 1.2212146e-08, 0.00015893648, -3.506652e-05, -9.288302e-06, 4.5798282e-07, 2.875361e-07, 1.7444851e-08};
endpackage
`endif
