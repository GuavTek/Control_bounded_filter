`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam N = 4;
	localparam real hf[0:1599] = {7.287086e-05, -5.8787242e-05, 9.878951e-06, -4.915542e-07, 4.4587272e-05, -5.429356e-05, 1.0070655e-05, -6.230468e-07, 1.8628934e-05, -4.949859e-05, 1.0156337e-05, -7.481968e-07, -4.871819e-06, -4.4475535e-05, 1.0137675e-05, -8.6520987e-07, -2.5819232e-05, -3.9297345e-05, 1.0017847e-05, -9.724776e-07, -4.4153745e-05, -3.4035686e-05, 9.801415e-06, -1.068598e-06, -5.9851103e-05, -2.875996e-05, 9.494201e-06, -1.1523917e-06, -7.2921e-05, -2.3536437e-05, 9.103138e-06, -1.2229137e-06, -8.340531e-05, -1.8427434e-05, 8.636113e-06, -1.2794591e-06, -9.137594e-05, -1.3490627e-05, 8.10181e-06, -1.3215655e-06, -9.6932316e-05, -8.778441e-06, 7.5095327e-06, -1.3490114e-06, -0.00010019868, -4.3375626e-06, 6.86904e-06, -1.3618096e-06, -0.0001013211, -2.0855683e-07, 6.1903725e-06, -1.3601974e-06, -0.00010046431, 3.5744063e-06, 5.4836883e-06, -1.3446232e-06, -9.780854e-05, 6.9837133e-06, 4.759102e-06, -1.315731e-06, -9.3546114e-05, 9.998366e-06, 4.0265327e-06, -1.2743407e-06, -8.787825e-05, 1.2603938e-05, 3.2955654e-06, -1.2214283e-06, -8.1011756e-05, 1.479243e-05, 2.575319e-06, -1.1581031e-06, -7.315585e-05, 1.6562048e-05, 1.8743342e-06, -1.0855845e-06, -6.451918e-05, 1.7916891e-05, 1.200472e-06, -1.0051772e-06, -5.530696e-05, 1.8866573e-05, 5.6082973e-07, -9.182474e-07, -4.571828e-05, 1.942578e-05, -3.8326775e-08, -8.261983e-07, -3.594373e-05, 1.9613777e-05, -5.916148e-07, -7.304462e-07, -2.6163243e-05, 1.9453879e-05, -1.0945699e-06, -6.3239787e-07, -1.6544187e-05, 1.897288e-05, -1.5436647e-06, -5.334293e-07, -7.2397925e-06, 1.8200471e-05, -1.936312e-06, -4.348651e-07, 1.6121634e-06, 1.7168648e-05, -2.2708537e-06, -3.3796107e-07, 9.8903465e-06, 1.591111e-05, -2.5465351e-06, -2.4388777e-07, 1.7490578e-05, 1.44626765e-05, -2.7634674e-06, -1.5371661e-07, 2.432625e-05, 1.2858717e-05, -2.9225778e-06, -6.840838e-08, 3.032846e-05, 1.1134606e-05, -3.0255508e-06, 1.1195987e-08, 3.5445886e-05, 9.32521e-06, -3.0747608e-06, 8.438222e-08, 3.9644416e-05, 7.4644113e-06, -3.073197e-06, 1.5056705e-07, 4.2906533e-05, 5.5846767e-06, -3.0243841e-06, 2.0930023e-07, 4.5230525e-05, 3.7166722e-06, -2.9322994e-06, 2.6026433e-07, 4.6629484e-05, 1.8889268e-06, -2.8012864e-06, 3.0327243e-07, 4.713018e-05, 1.2755018e-07, -2.6359698e-06, 3.3826362e-07, 4.6771773e-05, -1.5439988e-06, -2.441169e-06, 3.6529704e-07, 4.560446e-05, -3.1050874e-06, -2.221816e-06, 3.8454405e-07, 4.3688015e-05, -4.538034e-06, -1.9828747e-06, 3.962791e-07, 4.1090294e-05, -5.8281776e-06, -1.7292665e-06, 4.0086948e-07, 3.7885733e-05, -6.963904e-06, -1.4657992e-06, 3.987642e-07, 3.4153807e-05, -7.936622e-06, -1.1971035e-06, 3.9048206e-07, 2.997755e-05, -8.740692e-06, -9.275761e-07, 3.7659942e-07, 2.5442092e-05, -9.373324e-06, -6.613292e-07, 3.5773758e-07, 2.0633279e-05, -9.83444e-06, -4.0214903e-07, 3.3455055e-07, 1.5636351e-05, -1.012649e-05, -1.5346086e-07, 3.0771253e-07, 1.0534734e-05, -1.0254266e-05, 8.1697415e-08, 2.7790625e-07, 5.4089137e-06, -1.0224679e-05, 3.0069407e-07, 2.458118e-07, 3.3544268e-07, -1.0046516e-05, 5.0131484e-07, 2.1209594e-07, -4.61394e-06, -9.730204e-06, 6.817672e-07, 1.7740277e-07, -9.373064e-06, -9.287546e-06, 8.406773e-07, 1.4234493e-07, -1.38819505e-05, -8.731468e-06, 9.770812e-07, 1.0749628e-07, -1.8087312e-05, -8.075762e-06, 1.0904104e-06, 7.3385365e-08, -2.1942918e-05, -7.3348288e-06, 1.1804716e-06, 4.0490345e-08, -2.5409843e-05, -6.5234417e-06, 1.2474236e-06, 9.234943e-09, -2.8456589e-05, -5.6565113e-06, 1.2917486e-06, -2.0014351e-08, -3.10591e-05, -4.7488675e-06, 1.3142222e-06, -4.694994e-08, -3.3200675e-05, -3.8150583e-06, 1.3158806e-06, -7.1323676e-08, -3.487178e-05, -2.869166e-06, 1.2979862e-06, -9.2946365e-08, -3.6069767e-05, -1.9246431e-06, 1.2619923e-06, -1.1168634e-07, -3.679852e-05, -9.94168e-07, 1.2095084e-06, -1.2746713e-07, -3.706805e-05, -8.952218e-08, 1.1422648e-06, -1.4026436e-07, -3.6894016e-05, 7.7851183e-07, 1.0620789e-06, -1.5010205e-07, -3.6297188e-05, 1.6002319e-06, 9.708227e-07, -1.5704833e-07, -3.5302914e-05, 2.3670768e-06, 8.7039245e-07, -1.6121074e-07, -3.3940523e-05, 3.0716678e-06, 7.626796e-07, -1.6273118e-07, -3.2242737e-05, 3.7078305e-06, 6.4954537e-07, -1.6178082e-07, -3.0245052e-05, 4.2706006e-06, 5.327973e-07, -1.5855467e-07, -2.798516e-05, 4.7562125e-06, 4.141687e-07, -1.5326646e-07, -2.550233e-05, 5.162073e-06, 2.953012e-07, -1.4614345e-07, -2.2836846e-05, 5.486725e-06, 1.7772989e-07, -1.3742148e-07, -2.0029449e-05, 5.7297934e-06, 6.287174e-08, -1.273404e-07, -1.7120803e-05, 5.89193e-06, -4.7983598e-08, -1.16139674e-07, -1.4151011e-05, 5.974741e-06, -1.5368006e-07, -1.0405459e-07, -1.11591435e-05, 5.9807144e-06, -2.5319912e-07, -9.131275e-08, -8.1828275e-06, 5.9131403e-06, -3.456614e-07, -7.8131116e-08, -5.257859e-06, 5.776027e-06, -4.303262e-07, -6.471355e-08, -2.417871e-06, 5.574015e-06, -5.065893e-07, -5.1248783e-08, 3.059652e-07, 5.3122903e-06, -5.7397915e-07, -3.7908983e-08, 2.8851878e-06, 4.996495e-06, -6.321518e-07, -2.4848674e-08, 5.2942532e-06, 4.632646e-06, -6.8088457e-07, -1.2204211e-08, 7.5107014e-06, 4.2270444e-06, -7.200691e-07, -9.3608093e-11, 9.515276e-06, 3.786199e-06, -7.4970404e-07, 1.1383223e-08, 1.1292012e-05, 3.316743e-06, -7.698865e-07, 2.2143913e-08, 1.2828272e-05, 2.8253605e-06, -7.8080444e-07, 3.2122788e-08, 1.4114763e-05, 2.3187154e-06, -7.827279e-07, 4.1269775e-08, 1.5145501e-05, 1.8033815e-06, -7.760013e-07, 4.9549147e-08, 1.5917754e-05, 1.285782e-06, -7.6103515e-07, 5.6938124e-08, 1.6431952e-05, 7.721297e-07, -7.382988e-07, 6.342538e-08, 1.6691567e-05, 2.6837301e-07, -7.0831277e-07, 6.9009566e-08, 1.6702967e-05, -2.1985295e-07, -6.7164206e-07, 7.369777e-08, 1.6475253e-05, -6.8727115e-07, -6.288897e-07, 7.750413e-08, 1.6020062e-05, -1.1290025e-06, -5.8069054e-07, 8.044844e-08, 1.5351368e-05, -1.5406013e-06, -5.277055e-07, 8.255493e-08, 1.4485251e-05, -1.9180857e-06, -4.706163e-07, 8.3851184e-08, 1.34396605e-05, -2.257964e-06, -4.1012038e-07, 8.436723e-08, 1.2234164e-05, -2.5572567e-06, -3.4692584e-07, 8.413474e-08, 1.0889689e-05, -2.813512e-06, -2.8174685e-07, 8.318651e-08, 9.428253e-06, -3.0248202e-06, -2.152991e-07, 8.155599e-08, 7.872692e-06, -3.1898194e-06, -1.4829513e-07, 7.927712e-08, 6.246384e-06, -3.3077006e-06, -8.143986e-08, 7.638421e-08, 4.5729757e-06, -3.3782053e-06, -1.5425996e-08, 7.291201e-08, 2.8761049e-06, -3.4016196e-06, 4.9070643e-08, 6.8895915e-08, 1.1791337e-06, -3.3787633e-06, 1.113959e-07, 6.437221e-08, -4.951165e-07, -3.3109748e-06, 1.7092209e-07, 5.937845e-08, -2.1246185e-06, -3.2000908e-06, 2.27053e-07, 5.3953855e-08, -3.688383e-06, -3.0484216e-06, 2.7922886e-07, 4.8139682e-08, -5.1666875e-06, -2.8587215e-06, 3.2693134e-07, 4.197966e-08, -6.541292e-06, -2.6341559e-06, 3.6968865e-07, 3.5520323e-08, -7.795632e-06, -2.3782625e-06, 4.0708034e-07, 2.8811307e-08, -8.914999e-06, -2.0949096e-06, 4.3874215e-07, 2.1905556e-08, -9.886688e-06, -1.7882513e-06, 4.6437037e-07, 1.4859423e-08, -1.0700135e-05, -1.4626769e-06, 4.83726e-07, 7.732637e-09, -1.1347019e-05, -1.12276e-06, 4.9663856e-07, 5.8815736e-10, -1.18213375e-05, -7.7320317e-07, 5.0300883e-07, -6.508126e-09, -1.2119463e-05, -4.1878243e-07, 5.028118e-07, -1.3487834e-08, -1.2240161e-05, -6.428836e-08, 4.960982e-07, -2.0280675e-08, -1.2184583e-05, 2.8553202e-07, 4.829952e-07, -2.6815165e-08, -1.1956232e-05, 6.260341e-07, 4.6370664e-07, -3.3019468e-08, -1.1560896e-05, 9.527335e-07, 4.3851216e-07, -3.882234e-08, -1.1006553e-05, 1.2613631e-06, 4.0776496e-07, -4.415418e-08, -1.0303248e-05, 1.5479269e-06, 3.718889e-07, -4.8948127e-08, -9.462946e-06, 1.808752e-06, 3.3137448e-07, -5.3141235e-08, -8.499358e-06, 2.0405364e-06, 2.8677363e-07, -5.667563e-08, -7.4277445e-06, 2.2403922e-06, 2.3869364e-07, -5.949969e-08, -6.2646986e-06, 2.405884e-06, 1.8778994e-07, -6.156916e-08, -5.02791e-06, 2.535062e-06, 1.3475827e-07, -6.284822e-08, -3.7359175e-06, 2.6264875e-06, 8.032572e-08, -6.331048e-08, -2.407847e-06, 2.6792532e-06, 2.5241325e-08, -6.293977e-08, -1.0631422e-06, 2.6929952e-06, -2.973403e-08, -6.1730894e-08, 2.7870774e-07, 2.6678983e-06, -8.383808e-08, -5.9690166e-08, 1.5984429e-06, 2.604693e-06, -1.3631791e-07, -5.6835717e-08, 2.877303e-06, 2.504645e-06, -1.8644081e-07, -5.31977e-08, 4.0972905e-06, 2.3695372e-06, -2.3350502e-07, -4.8818187e-08, 5.241424e-06, 2.201644e-06, -2.768502e-07, -4.3750916e-08, 6.293974e-06, 2.003698e-06, -3.1586748e-07, -3.8060783e-08, 7.240686e-06, 1.7788506e-06, -3.5000897e-07, -3.1823127e-08, 8.068974e-06, 1.5306255e-06, -3.787964e-07, -2.5122805e-08, 8.768098e-06, 1.2628669e-06, -4.0182863e-07, -1.8053063e-08, 9.329308e-06, 9.796831e-07, -4.1878857e-07, -1.0714238e-08, 9.7459615e-06, 6.8538486e-07, -4.294484e-07, -3.2122875e-09, 1.00136085e-05, 3.8442158e-07, -4.3367362e-07, 4.342815e-09, 1.0130045e-05, 8.131475e-08, -4.3142572e-07, 1.1838793e-08, 1.0095331e-05, -2.1940977e-07, -4.2276335e-07, 1.9162858e-08, 9.911778e-06, -5.1328976e-07, -4.0784184e-07, 2.6203557e-08, 9.583898e-06, -7.9599374e-07, -3.8691135e-07, 3.2852615e-08, 9.118322e-06, -1.0633861e-06, -3.6031344e-07, 3.9006775e-08, 8.523687e-06, -1.3115896e-06, -3.284759e-07, 4.4569585e-08, 7.810492e-06, -1.5370432e-06, -2.9190656e-07, 4.9453064e-08, 6.9909283e-06, -1.736556e-06, -2.5118555e-07, 5.357929e-08, 6.0786765e-06, -1.9073545e-06, -2.0695623e-07, 5.6881795e-08, 5.088694e-06, -2.0471236e-06, -1.5991526e-07, 5.9306817e-08, 4.0369714e-06, -2.1540413e-06, -1.10801665e-07, 6.081431e-08, 2.940284e-06, -2.226804e-06, -6.0385105e-08, 6.1378735e-08, 1.8159244e-06, -2.2646443e-06, -9.453677e-09, 6.098965e-08, 6.814323e-07, -2.2673412e-06, 4.1198653e-08, 5.965196e-08, -4.4567847e-07, -2.2352199e-06, 9.078478e-08, 5.7385993e-08, -1.5481921e-06, -2.1691449e-06, 1.3853708e-07, 5.4227225e-08, -2.6094563e-06, -2.0705022e-06, 1.837197e-07, 5.0225804e-08, -3.613637e-06, -1.9411752e-06, 2.2564049e-07, 4.5445777e-08, -4.5459606e-06, -1.7835122e-06, 2.6366203e-07, 3.996408e-08, -5.3929343e-06, -1.6002856e-06, 2.9721187e-07, 3.3869295e-08, -6.1425494e-06, -1.3946459e-06, 3.2579172e-07, 2.7260219e-08, -6.784455e-06, -1.1700685e-06, 3.4898537e-07, 2.0244205e-08, -7.3101073e-06, -9.3029627e-07, 3.6646517e-07, 1.2935382e-08, -7.71289e-06, -6.7927806e-07, 3.779972e-07, 5.452746e-09, -7.988196e-06, -4.2110346e-07, 3.834447e-07, -2.0818551e-09, -8.133487e-06, -1.5993656e-07, 3.8277003e-07, -9.54578e-09, -8.148312e-06, 1.0005182e-07, 3.7603476e-07, -1.6817676e-08, -8.034292e-06, 3.547514e-07, 3.6339839e-07, -2.3779537e-08, -7.795073e-06, 6.0017817e-07, 3.4511513e-07, -3.031871e-08, -7.436249e-06, 8.3253803e-07, 3.2152934e-07, -3.6329812e-08, -6.9652524e-06, 1.0482864e-06, 2.9306935e-07, -4.1716515e-08, -6.3912134e-06, 1.2441839e-06, 2.6023991e-07, -4.639318e-08, -5.7247953e-06, 1.4173459e-06, 2.2361343e-07, -5.0286296e-08, -4.978004e-06, 1.5652864e-06, 1.8382e-07, -5.333572e-08, -4.1639837e-06, 1.6859557e-06, 1.415367e-07, -5.5495672e-08, -3.296786e-06, 1.7777684e-06, 9.747591e-08, -5.6735466e-08, -2.3911352e-06, 1.839626e-06, 5.237329e-08, -5.704002e-08, -1.4621808e-06, 1.8709294e-06, 6.9753345e-09, -5.6410023e-08, -5.252445e-07, 1.8715843e-06, -3.797317e-08, -5.486192e-08, 4.0442933e-07, 1.8419975e-06, -8.1741575e-08, -5.2427524e-08, 1.3119233e-06, 1.7830645e-06, -1.2362547e-07, -4.9153424e-08, 2.1828857e-06, 1.6961503e-06, -1.6295832e-07, -4.510013e-08, 3.0037595e-06, 1.5830615e-06, -1.9912227e-07, -4.034095e-08, 3.761994e-06, 1.4460114e-06, -2.3155815e-07, -3.496069e-08, 4.4462395e-06, 1.2875796e-06, -2.5977437e-07, -2.9054103e-08, 5.046516e-06, 1.1106645e-06, -2.833546e-07, -2.2724246e-08, 5.554364e-06, 9.184314e-07, -3.019641e-07, -1.6080625e-08, 5.9629606e-06, 7.1425774e-07, -3.1535458e-07, -9.237292e-09, 6.2672134e-06, 5.0167347e-07, -3.2336766e-07, -2.3108406e-09, 6.4638202e-06, 2.8430094e-07, -3.2593664e-07, 4.581613e-09, 6.5512995e-06, 6.579329e-08, -3.230867e-07, 1.1324453e-08, 6.5299932e-06, -1.5022708e-07, -3.1493366e-07, 1.780555e-08, 6.402033e-06, -3.6022854e-07, -3.0168098e-07, 2.3918169e-08, 6.1712813e-06, -5.608283e-07, -2.8361552e-07, 2.9562768e-08, 5.8432447e-06, -7.488472e-07, -2.6110166e-07, 3.4648664e-08, 5.4249563e-06, -9.213605e-07, -2.3457451e-07, 3.909554e-08, 4.9248392e-06, -1.0757435e-06, -2.0453152e-07, 4.283472e-08, 4.3525456e-06, -1.2097124e-06, -1.7152338e-07, 4.5810296e-08, 3.7187763e-06, -1.3213573e-06, -1.3614421e-07, 4.7979956e-08, 3.0350884e-06, -1.4091703e-06, -9.9020696e-08, 4.931562e-08, 2.3136881e-06, -1.4720649e-06, -6.080123e-08, 4.9803777e-08, 1.5672164e-06, -1.5093893e-06, -2.2144457e-08, 4.9445603e-08, 8.0853044e-07, -1.5209308e-06, 1.6292034e-08, 4.8256787e-08, 5.048438e-08, -1.5069137e-06, 5.3862973e-08, 4.6267136e-08, -6.942873e-07, -1.4679891e-06, 8.994629e-08, 4.351991e-08, -1.4135792e-06, -1.4052187e-06, 1.239535e-07, 4.0070937e-08, -2.0958141e-06, -1.3200496e-06, 1.5533936e-07, 3.5987515e-08, -2.7302292e-06, -1.2142855e-06, 1.8361071e-07, 3.134713e-08, -3.3070455e-06, -1.0900502e-06, 2.0833424e-07, 2.6235998e-08, -3.8176167e-06, -9.497469e-07, 2.2914318e-07, 2.074747e-08, -4.25456e-06, -7.960133e-07, 2.4574277e-07, 1.498033e-08, -4.611859e-06, -6.316731e-07, 2.579144e-07, 9.037017e-09, -4.8849456e-06, -4.59685e-07, 2.6551828e-07, 3.0217988e-09, -5.070755e-06, -2.8309026e-07, 2.6849494e-07, -2.9610716e-09, -5.1677503e-06, -1.0495927e-07, 2.6686502e-07, -8.8091685e-09, -5.175928e-06, 7.1661205e-08, 2.6072794e-07, -1.4423664e-08, -5.096791e-06, 2.4379997e-07, 2.5025906e-07, -1.9711011e-08, -4.933298e-06, 4.0861116e-07, 2.357056e-07, -2.4584516e-08, -4.6897903e-06, 5.6342105e-07, 2.1738133e-07, -2.8965768e-08, -4.371893e-06, 7.057713e-07, 1.9566026e-07, -3.278592e-08, -3.986399e-06, 8.334579e-07, 1.7096927e-07, -3.598676e-08, -3.5411329e-06, 9.445648e-07, 1.4377996e-07, -3.8521616e-08, -3.044798e-06, 1.0374927e-06, 1.14599835e-07, -4.0356017e-08, -2.5068143e-06, 1.110981e-06, 8.396295e-08, -4.1468148e-08, -1.9371435e-06, 1.1641246e-06, 5.2420283e-08, -4.184907e-08, -1.3461091e-06, 1.1963836e-06, 2.0529871e-08, -4.1502705e-08, -7.4421206e-07, 1.207586e-06, -1.1152979e-08, -4.0445617e-08, -1.4194762e-07, 1.1979262e-06, -4.2085322e-08, -3.8706524e-08, 4.503754e-07, 1.1679538e-06, -7.174584e-08, -3.632567e-08, 1.0228092e-06, 1.1185592e-06, -9.96436e-08, -3.3353935e-08, 1.5659322e-06, 1.0509527e-06, -1.2532617e-07, -2.9851815e-08, 2.0710022e-06, 9.666373e-07, -1.4838687e-07, -2.588821e-08, 2.530096e-06, 8.673787e-07, -1.6847126e-07, -2.1539114e-08, 2.936231e-06, 7.551691e-07, -1.8528245e-07, -1.6886169e-08, 3.2834703e-06, 6.321896e-07, -1.9858537e-07, -1.2015151e-08, 3.5670057e-06, 5.0076886e-07, -2.0821e-07, -7.0143993e-09, 3.7832217e-06, 3.6333975e-07, -2.1405326e-07, -1.973225e-09, 3.9297356e-06, 2.2239543e-07, -2.1607977e-07, 3.0196787e-09, 4.0054183e-06, 8.044476e-08, -2.1432136e-07, 7.8777935e-09, 4.0103887e-06, -6.003169e-08, -2.0887549e-07, 1.2518272e-08, 3.9459906e-06, -1.9662446e-07, -1.9990242e-07, 1.6863346e-08, 3.814746e-06, -3.2703608e-07, -1.8762141e-07, 2.0841632e-08, 3.62029e-06, -4.4911923e-07, -1.7230593e-07, 2.4389289e-08, 3.3672864e-06, -5.6091164e-07, -1.5427791e-07, 2.7451046e-08, 3.061327e-06, -6.6066724e-07, -1.3390131e-07, 2.998105e-08, 2.7088174e-06, -7.4688273e-07, -1.1157499e-07, 3.194353e-08, 2.316849e-06, -8.1831985e-07, -8.7725184e-08, 3.3313288e-08, 1.8930629e-06, -8.740222e-07, -6.279742e-08, 3.4075985e-08, 1.445505e-06, -9.133268e-07, -3.7248412e-08, 3.4228226e-08, 9.824778e-07, -9.3587084e-07, -1.1537805e-08, 3.377745e-08, 5.1239016e-07, -9.415922e-07, 1.3880017e-08, 3.2741635e-08, 4.3607365e-08, -9.3072543e-07, 3.8563854e-08, 3.114882e-08, -4.1569484e-07, -9.0379194e-07, 6.2093264e-08, 2.9036443e-08, -8.576703e-07, -8.6158565e-07, 8.407566e-08, 2.645054e-08, -1.2749341e-06, -8.0515395e-07, 1.0415275e-07, 2.3444777e-08, -1.6606838e-06, -7.3577473e-07, 1.2200634e-07, 2.0079387e-08, -2.008808e-06, -6.549293e-07, 1.3736324e-07, 1.6419994e-08, -2.313981e-06, -5.642726e-07, 1.4999935e-07, 1.253635e-08, -2.5717404e-06, -4.6560066e-07, 1.5974277e-07, 8.501036e-09, -2.7785513e-06, -3.6081622e-07, 1.6647596e-07, 4.3881223e-09, -2.9318487e-06, -2.5189294e-07, 1.7013686e-07, 2.7182026e-10, -3.0300648e-06, -1.408393e-07, 1.7071899e-07, -3.7748396e-09, -3.0726371e-06, -2.9662125e-08, 1.6827067e-07, -7.681292e-09, -3.059999e-06, 7.966887e-08, 1.6289313e-07, -1.1380659e-08, -2.9935522e-06, 1.8525542e-07, 1.5473775e-07, -1.4810878e-08, -2.8756228e-06, 2.85303e-07, 1.4400256e-07, -1.7915738e-08, -2.7094025e-06, 3.781509e-07, 1.3092775e-07, -2.0645784e-08, -2.4988733e-06, 4.6229908e-07, 1.15790776e-07, -2.2959087e-08, -2.2487227e-06, 5.364319e-07, 9.890064e-08, -2.4821876e-08, -1.9642457e-06, 5.994381e-07, 8.059186e-08, -2.6209003e-08, -1.6512383e-06, 6.504266e-07, 6.121798e-08, -2.7104246e-08, -1.3158843e-06, 6.887381e-07, 4.1144975e-08, -2.7500455e-08, -9.646378e-07, 7.139527e-07, 2.0744425e-08, -2.7399526e-08, -6.041021e-07, 7.2589245e-07, 3.8679684e-10, -2.6812215e-08, -2.4090937e-07, 7.2462007e-07, -1.9565183e-08, -2.5757792e-08, 1.1839895e-07, 7.104332e-07, -3.8762884e-08, -2.4263555e-08, 4.6748684e-07, 6.8385447e-07, -5.6877756e-08, -2.2364201e-08, 8.0033317e-07, 6.4561766e-07, -7.360687e-08, -2.010108e-08, 1.1113331e-06, 5.966508e-07, -8.8677865e-08, -1.7521334e-08, 1.3953901e-06, 5.380553e-07, -1.0185329e-07, -1.467695e-08, 1.647997e-06, 4.7108333e-07, -1.1293422e-07, -1.1623749e-08, 1.8653052e-06, 3.9711185e-07, -1.2176314e-07, -8.420307e-09, 2.0441805e-06, 3.176159e-07, -1.2822596e-07, -5.126859e-09, 2.1822443e-06, 2.3413997e-07, -1.3225338e-07, -1.8041821e-09, 2.2779022e-06, 1.482688e-07, -1.3382113e-07, 1.4875061e-09, 2.3303558e-06, 6.159819e-08, -1.3294975e-07, 4.6896247e-09, 2.3396015e-06, -2.4294005e-08, -1.297033e-07, 7.746255e-09, 2.3064142e-06, -1.0787598e-07, -1.2418735e-07, 1.0605108e-08, 2.232318e-06, -1.8768866e-07, -1.1654643e-07, 1.3218395e-08, 2.1195422e-06, -2.6237063e-07, -1.0696059e-07, 1.5543622e-08, 1.9709687e-06, -3.306808e-07, -9.564151e-08, 1.7544254e-08, 1.7900653e-06, -3.915184e-07, -8.28281e-08, 1.919028e-08, 1.580811e-06, -4.439402e-07, -6.878167e-08, 2.0458632e-08, 1.3476148e-06, -4.871744e-07, -5.378075e-08, 2.1333484e-08, 1.0952259e-06, -5.206313e-07, -3.8115775e-08, 2.1806413e-08, 8.2864136e-07, -5.4391023e-07, -2.2083572e-08, 2.1876408e-08, 5.530107e-07, -5.5680323e-07, -5.981872e-09, 2.1549772e-08, 2.7353886e-07, -5.59295e-07, 9.896111e-09, 2.0839867e-08, -4.6088555e-09, -5.5155925e-07, 2.5266898e-08, 1.9766752e-08, -2.7640007e-07, -5.339519e-07, 3.9861717e-08, 1.8356696e-08, -5.370239e-07, -5.0700106e-07, 5.34311e-08, 1.6641593e-08, -7.8197394e-07, -4.7139395e-07, 6.574904e-08, 1.4658282e-08, -1.0071241e-06, -4.279612e-07, 7.661667e-08, 1.2447789e-08, -1.2087955e-06, -3.776591e-07, 8.586535e-08, 1.0054508e-08, -1.3838153e-06, -3.2154944e-07, 9.335917e-08, 7.525337e-09, -1.5295632e-06, -2.607783e-07, 9.89968e-08, 4.9087725e-09, -1.6440082e-06, -1.965535e-07, 1.0271268e-07, 2.254007e-09, -1.7257341e-06, -1.3012112e-07, 1.0447754e-07, -3.8998144e-10, -1.7739527e-06, -6.274226e-08, 1.04298245e-07, -2.9753164e-09, -1.7885046e-06, 4.330382e-09, 1.02216966e-07, -5.456074e-09, -1.7698507e-06, 6.9875206e-08, 9.830977e-08, -7.789084e-09, -1.7190498e-06, 1.3272341e-07, 9.268457e-08, -9.934666e-09, -1.6377279e-06, 1.9177934e-07, 8.5478554e-08, -1.1857293e-08, -1.5280367e-06, 2.4603898e-07, 7.685514e-08, -1.3526154e-08, -1.3926033e-06, 2.946067e-07, 6.700044e-08, -1.4915646e-08, -1.2344728e-06, 3.367093e-07, 5.611951e-08, -1.6005728e-08, -1.0570435e-06, 3.7170793e-07, 4.4432163e-08, -1.6782202e-08, -8.6399785e-07, 3.9910697e-07, 3.216871e-08, -1.7236857e-08, -6.592286e-07, 4.1856052e-07, 1.9565531e-08, -1.7367515e-08, -4.4676355e-07, 4.298755e-07, 6.860638e-09, -1.7177953e-08, -2.3068839e-07, 4.3301253e-07, -5.7107257e-09, -1.6677738e-08, -1.5070663e-08, 4.280832e-07, -1.7920334e-08, -1.5881936e-08, 1.9611478e-07, 4.1534545e-07, -2.9551035e-08, -1.4810738e-08, 3.9905714e-07, 3.951957e-07, -4.0400522e-08, -1.3489006e-08, 5.9017634e-07, 3.6815896e-07, -5.028476e-08, -1.1945721e-08, 7.6618466e-07, 3.3487646e-07, -5.904103e-08, -1.0213382e-08, 9.241411e-07, 2.9609183e-07, -6.65305e-08, -8.32735e-09, 1.0614989e-06, 2.526352e-07, -7.264032e-08, -6.3251435e-09, 1.1761443e-06, 2.0540631e-07, -7.7285215e-08, -4.245711e-09, 1.2664277e-06, 1.5535645e-07, -8.040853e-08, -2.1286948e-09, 1.3311835e-06, 1.0347004e-07, -8.1982726e-08, -1.3687354e-11, 1.3697432e-06, 5.0745776e-08, -8.200933e-08, 2.0604924e-09, 1.3819372e-06, -1.8221163e-09, -8.051835e-08, 4.0564982e-09, 1.3680881e-06, -5.3262102e-08, -7.7567215e-08, 5.9391145e-09, 1.3289948e-06, -1.02642865e-07, -7.323918e-08, 7.675865e-09, 1.2659086e-06, -1.490897e-07, -6.764129e-08, 9.237559e-09, 1.1805009e-06, -1.9179964e-07, -6.0901975e-08, 1.059877e-08, 1.0748236e-06, -2.3005484e-07, -5.316828e-08, 1.1738228e-08, 9.5126364e-07, -2.6323423e-07, -4.460279e-08, 1.2639145e-08, 8.1249266e-07, -2.9082318e-07, -3.538035e-08, 1.3289432e-08, 6.6141126e-07, -3.1242087e-07, -2.568459e-08, 1.3681841e-08, 5.0109065e-07, -3.277456e-07, -1.5704387e-08, 1.3814012e-08, 3.3471267e-07, -3.3663764e-07, -5.6302643e-09, 1.3688421e-08, 1.6550823e-07, -3.3905994e-07, 4.349157e-09, 1.3312252e-08, -3.30363e-09, -3.350963e-07, 1.4050604e-08, 1.2697174e-08, -1.6857521e-07, -3.2494765e-07, 2.3299448e-08, 1.185905e-08, -3.2728738e-07, -3.0892596e-07, 3.1932764e-08, 1.0817563e-08, -4.7660322e-07, -2.8744637e-07, 3.980214e-08, 9.5957855e-09, -6.1391717e-07, -2.6101748e-07, 4.6776126e-08, 8.2196925e-09, -7.3689915e-07, -2.3023017e-07, 5.2742386e-08, 6.7176296e-09, -8.4353235e-07, -1.9574503e-07, 5.7609398e-08, 5.1197446e-09, -9.3214516e-07, -1.582787e-07, 6.1307766e-08, 3.4574015e-09, -1.0014351e-06, -1.18589526e-07, 6.37911e-08, 1.7625765e-09, -1.0504863e-06, -7.746273e-08, 6.503644e-08, 6.725737e-11, -1.0787792e-06, -3.5695177e-08, 6.504425e-08, -1.5971476e-09, -1.0861925e-06, 5.9195933e-09, 6.383797e-08, -3.2003802e-09, -1.0729974e-06, 4.6606097e-08, 6.146318e-08, -4.71387e-09, -1.039846e-06, 8.562099e-08, 5.7986306e-08, -6.1112333e-09, -9.877507e-07, 1.2226631e-07, 5.3493025e-08, -7.368719e-09, -9.1805936e-07, 1.5590163e-07, 4.8086324e-08, -8.465604e-09, -8.3242327e-07, 1.8595487e-07, 4.188425e-08, -9.384519e-09, -7.327606e-07, 2.1193176e-07, 3.501745e-08, -1.0111711e-08, -6.212158e-07, 2.334235e-07, 2.7626518e-08, -1.063723e-08, -5.0011477e-07, 2.5011283e-07, 1.985919e-08, -1.0955048e-08, -3.719184e-07, 2.6177827e-07, 1.1867465e-08, -1.1063101e-08, -2.3917374e-07, 2.682964e-07, 3.804716e-09, -1.0963248e-08, -1.04464995e-07, 2.6964236e-07, -4.1772044e-09, -1.0661176e-08, 2.9635752e-08, 2.6588856e-07, -1.193075e-08, -1.0166218e-08, 1.6061624e-07, 2.5720144e-07, -1.9315348e-08, -9.491121e-09, 2.8607002e-07, 2.4383664e-07, -2.6199896e-08, -8.65174e-09, 4.037395e-07, 2.2613264e-07, -3.2465014e-08, -7.6666975e-09, 5.115554e-07, 2.0450281e-07, -3.8005073e-08, -6.5569816e-09, 6.0767206e-07, 1.7942641e-07, -4.2729894e-08, -5.3455187e-09, 6.9049787e-07, 1.514384e-07, -4.6566157e-08, -4.0567096e-09, 7.5872026e-07, 1.211184e-07, -4.9458464e-08, -2.7159535e-09, 8.113254e-07, 8.907905e-08, -5.1370037e-08, -1.3491561e-09, 8.476114e-07, 5.5953972e-08, -5.228307e-08, 1.7758107e-11, 8.67196e-07, 2.2385537e-08, -5.2198736e-08, 1.3593294e-09, 8.700178e-07, -1.0987314e-08, -5.1136794e-08, 2.6510265e-09, 8.563315e-07, -4.354095e-08, -4.913491e-08, 3.869686e-09, 8.266975e-07, -7.467844e-08, -4.6247624e-08, 4.993918e-09, 7.819655e-07, -1.0384022e-07, -4.2545032e-08, 6.004474e-09, 7.23254e-07, -1.3051393e-07, -3.8111207e-08, 6.8845623e-09, 6.5192376e-07, -1.542431e-07, -3.3042365e-08, 7.620122e-09, 5.695482e-07, -1.7463472e-07, -2.744487e-08, 8.200034e-09, 4.7788023e-07, -1.9136547e-07, -2.1433065e-08, 8.616273e-09, 3.7881577e-07, -2.0418646e-07, -1.5126991e-08, 8.864005e-09, 2.7435595e-07, -2.1292666e-07, -8.6500505e-09, 8.941622e-09, 1.6656755e-07, -2.1749463e-07, -2.1266435e-09, 8.850711e-09, 5.7542994e-08, -2.1787885e-07, 4.3201727e-09, 8.595973e-09, -5.063926e-08, -2.1414651e-07, 1.05709566e-08, 8.185076e-09, -1.5595356e-07, -2.0644089e-07, 1.6512047e-08, 7.628464e-09, -2.5646406e-07, -1.9497725e-07, 2.2037586e-08, 6.9391133e-09, -3.5035956e-07, -1.8003763e-07, 2.7051358e-08, 6.132243e-09, -4.3598524e-07, -1.6196434e-07, 3.1468417e-08, 5.2249973e-09, -5.1187095e-07, -1.4115246e-07, 3.5216473e-08, 4.2360897e-09, -5.7675567e-07, -1.18041555e-07, 3.8237022e-08, 3.1854277e-09};
	localparam real hb[0:1599] = {0.00010331091, -6.290727e-05, 9.581136e-06, -3.55674e-07, 0.00013570288, -6.6583234e-05, 9.178779e-06, -2.1749241e-07, 0.00016980777, -6.974785e-05, 8.675139e-06, -7.919704e-08, 0.00020535395, -7.233806e-05, 8.075186e-06, 5.695462e-08, 0.00024203959, -7.429614e-05, 7.385588e-06, 1.8866992e-07, 0.00027953554, -7.557086e-05, 6.6146804e-06, 3.136591e-07, 0.00031748883, -7.6118435e-05, 5.7723946e-06, 4.2967545e-07, 0.0003555267, -7.590356e-05, 4.870164e-06, 5.3455665e-07, 0.00039326103, -7.4900236e-05, 3.9207953e-06, 6.2626606e-07, 0.00043029318, -7.3092575e-05, 2.938312e-06, 7.029337e-07, 0.00046621924, -7.047539e-05, 1.9377733e-06, 7.628952e-07, 0.0005006355, -6.705473e-05, 9.350631e-07, 8.0472853e-07, 0.00053314405, -6.284816e-05, -5.3339015e-08, 8.2728735e-07, 0.00056335883, -5.7884965e-05, -1.0106075e-06, 8.297307e-07, 0.00059091125, -5.2206127e-05, -1.9198358e-06, 8.115475e-07, 0.0006154561, -4.5864108e-05, -2.764312e-06, 7.7257647e-07, 0.00063667726, -3.8922466e-05, -3.5278015e-06, 7.1301986e-07, 0.00065429293, -3.1455278e-05, -4.1948315e-06, 6.33451e-07, 0.00066806097, -2.3546363e-05, -4.750972e-06, 5.348159e-07, 0.0006777832, -1.528835e-05, -5.1831103e-06, 4.1842753e-07, 0.0006833099, -6.7815367e-06, -5.479711e-06, 2.8595343e-07, 0.0006845431, 1.867369e-06, -5.631059e-06, 1.3939693e-07, 0.0006814395, 1.0546687e-05, -5.6294784e-06, -1.8928743e-08, 0.00067401247, 1.9141306e-05, -5.469526e-06, -1.8643242e-07, 0.0006623335, 2.7534334e-05, -5.148151e-06, -3.6028305e-07, 0.00064653275, 3.560883e-05, -4.664822e-06, -5.374531e-07, 0.0006267983, 4.324959e-05, -4.0216105e-06, -7.1476677e-07, 0.0006033752, 5.0344952e-05, -3.2232397e-06, -8.8895246e-07, 0.00057656283, 5.6788605e-05, -2.277083e-06, -1.0566979e-06, 0.00054671225, 6.248136e-05, -1.1931227e-06, -1.214708e-06, 0.00051422184, 6.7332876e-05, 1.614004e-08, -1.3597644e-06, 0.00047953275, 7.1263246e-05, 1.3358185e-06, -1.4887834e-06, 0.000443123, 7.4204516e-05, 2.748819e-06, -1.5988754e-06, 0.0004055014, 7.610202e-05, 4.236061e-06, -1.6874006e-06, 0.00036720056, 7.691555e-05, 5.7767384e-06, -1.7520224e-06, 0.00032876927, 7.662031e-05, 7.3486135e-06, -1.7907561e-06, 0.0002907648, 7.520766e-05, 8.9283485e-06, -1.802013e-06, 0.00025374457, 7.2685645e-05, 1.0491859e-05, -1.784638e-06, 0.00021825773, 6.907921e-05, 1.2014691e-05, -1.7379406e-06, 0.00018483678, 6.443017e-05, 1.3472414e-05, -1.6617174e-06, 0.00015398912, 5.8796966e-05, 1.4841024e-05, -1.5562678e-06, 0.00012618888, 5.2254083e-05, 1.6097343e-05, -1.422399e-06, 0.00010186911, 4.48912e-05, 1.7219427e-05, -1.2614238e-06, 8.141446e-05, 3.6812107e-05, 1.818694e-05, -1.0751481e-06, 6.515442e-05, 2.8133367e-05, 1.8981538e-05, -8.6584953e-07, 5.335733e-05, 1.8982726e-05, 1.95872e-05, -6.362474e-07, 4.6225225e-05, 9.497333e-06, 1.9990544e-05, -3.894638e-07, 4.388964e-05, -1.782465e-07, 2.0181104e-05, -1.289767e-07, 4.640839e-05, -9.894159e-06, 2.015155e-05, 1.4143376e-07, 5.376352e-05, -1.9497527e-05, 1.9897874e-05, 4.1774595e-07, 6.586037e-05, -2.8834798e-05, 1.941952e-05, 6.957625e-07, 8.252781e-05, -3.775415e-05, 1.871945e-05, 9.711804e-07, 0.000103519764, -4.610791e-05, 1.7804161e-05, 1.239664e-06, 0.00012851782, -5.3754946e-05, 1.6683642e-05, 1.4969203e-06, 0.00015713515, -6.056299e-05, 1.5371268e-05, 1.7387738e-06, 0.00018892145, -6.6410874e-05, 1.3883635e-05, 1.9612412e-06, 0.00022336903, -7.1190596e-05, 1.2240336e-05, 2.1606031e-06, 0.0002599199, -7.4809235e-05, 1.04636965e-05, 2.3334724e-06, 0.00029797378, -7.71906e-05, 8.578441e-06, 2.476858e-06, 0.00033689666, -7.827672e-05, 6.611327e-06, 2.5882212e-06, 0.00037603045, -7.8028956e-05, 4.590736e-06, 2.6655257e-06, 0.00041470275, -7.642892e-05, 2.546232e-06, 2.7072797e-06, 0.0004522371, -7.3479e-05, 5.0809336e-07, 2.7125668e-06, 0.0004879635, -6.920259e-05, -1.4931725e-06, 2.6810694e-06, 0.0005212289, -6.3644e-05, -3.427324e-06, 2.6130808e-06, 0.0005514075, -5.6867975e-05, -5.2648816e-06, 2.5095057e-06, 0.0005779109, -4.895895e-05, -6.977618e-06, 2.3718505e-06, 0.0006001976, -4.0019935e-05, -8.539031e-06, 2.2022045e-06, 0.0006177818, -3.0171077e-05, -9.924795e-06, 2.0032069e-06, 0.00063024205, -1.9547972e-05, -1.1113176e-05, 1.7780077e-06, 0.0006372278, -8.299684e-06, -1.2085411e-05, 1.5302163e-06, 0.0006384661, 3.413466e-06, -1.2826043e-05, 1.2638432e-06, 0.0006337666, 1.542231e-05, -1.3323196e-05, 9.832337e-07, 0.000623025, 2.7551416e-05, -1.35688e-05, 6.9299455e-07, 0.0006062258, 3.962177e-05, -1.3558749e-05, 3.9791686e-07, 0.0005834434, 5.1453575e-05, -1.3293e-05, 1.02893665e-07, 0.0005548416, 6.286905e-05, -1.2775595e-05, -1.8716368e-07, 0.0005206722, 7.369521e-05, -1.2014624e-05, -4.6741047e-07, 0.0004812714, 8.3766674e-05, -1.1022117e-05, -7.331528e-07, 0.00043705595, 9.2928225e-05, -9.813865e-06, -9.799294e-07, 0.00038851702, 0.000101037345, -8.409186e-06, -1.20359e-06, 0.00033621336, 0.00010796651, -6.8306213e-06, -1.4003688e-06, 0.00028076337, 0.000113605274, -5.1035845e-06, -1.5669501e-06, 0.00022283595, 0.000117862044, -3.2559547e-06, -1.7005287e-06, 0.00016314084, 0.00012066564, -1.317631e-06, -1.7988592e-06, 0.00010241794, 0.00012196647, 6.799508e-07, -1.8602972e-06, 4.14264e-05, 0.00012173738, 2.7043286e-06, -1.8838289e-06, -1.9066772e-05, 0.000119974175, 4.722542e-06, -1.8690909e-06, -7.8298246e-05, 0.00011669572, 6.701672e-06, -1.8163773e-06, -0.00013551986, 0.000111943744, 8.609379e-06, -1.726637e-06, -0.0001900099, 0.00010578219, 1.0414434e-05, -1.6014574e-06, -0.000241084, 9.829629e-05, 1.2087232e-05, -1.4430381e-06, -0.00028810545, 8.959126e-05, 1.3600281e-05, -1.2541544e-06, -0.00033049483, 7.9790676e-05, 1.4928651e-05, -1.038109e-06, -0.00036773874, 6.903455e-05, 1.6050386e-05, -7.9867584e-07, -0.00039939737, 5.7477137e-05, 1.6946862e-05, -5.400348e-07, -0.00042511115, 4.5284574e-05, 1.7603095e-05, -2.666995e-07, -0.00044460606, 3.2632237e-05, 1.800799e-05, 1.6560573e-08, -0.00045769743, 1.9702016e-05, 1.8154506e-05, 3.0480268e-07, -0.00046429262, 6.679471e-06, 1.8039782e-05, 5.929965e-07, -0.00046439207, -6.249064e-06, 1.7665172e-05, 8.7611113e-07, -0.00045808902, -1.8899387e-05, 1.703622e-05, 1.149202e-06, -0.00044556762, -3.109229e-05, 1.6162558e-05, 1.4074968e-06, -0.00042709988, -4.2656346e-05, 1.5057738e-05, 1.6464774e-06, -0.00040304093, -5.3430525e-05, 1.3739011e-05, 1.8619577e-06, -0.0003738234, -6.3266685e-05, 1.2227024e-05, 2.050156e-06, -0.0003399502, -7.203182e-05, 1.0545476e-05, 2.2077593e-06, -0.0003019866, -7.961005e-05, 8.720718e-06, 2.33198e-06, -0.0002605512, -8.590433e-05, 6.7813157e-06, 2.4206036e-06, -0.00021630601, -9.083787e-05, 4.7575686e-06, 2.4720243e-06, -0.00016994624, -9.4355215e-05, 2.6810094e-06, 2.4852734e-06, -0.0001221893, -9.642295e-05, 5.838809e-07, 2.460033e-06, -7.3763695e-05, -9.7030046e-05, -1.5013957e-06, 2.396641e-06, -2.5397858e-05, -9.618793e-05, -3.5427522e-06, 2.2960826e-06, 2.2191041e-05, -9.393005e-05, -5.5089977e-06, 2.1599722e-06, 6.830793e-05, -9.031122e-05, -7.3703245e-06, 1.9905233e-06, 0.000112290254, -8.540655e-05, -9.098789e-06, 1.7905091e-06, 0.00015351785, -7.931006e-05, -1.0668757e-05, 1.5632132e-06, 0.0001914219, -7.213307e-05, -1.20573095e-05, 1.3123703e-06, 0.00022549325, -6.4002204e-05, -1.3244605e-05, 1.0421014e-06, 0.00025528937, -5.5057284e-05, -1.4214173e-05, 7.568419e-07, 0.0002804405, -4.5448956e-05, -1.495317e-05, 4.6126368e-07, 0.00030065438, -3.5336187e-05, -1.5452555e-05, 1.6019447e-07, 0.00031571978, -2.4883631e-05, -1.5707217e-05, -1.414653e-07, 0.00032550868, -1.4258976e-05, -1.5716014e-05, -4.3882665e-07, 0.00032997705, -3.6302097e-06, -1.548177e-05, -7.2709526e-07, 0.0003291644, 6.8370555e-06, -1.5011187e-05, -1.001653e-06, 0.00032319195, 1.6982198e-05, -1.4314705e-05, -1.2581353e-06, 0.0003122594, 2.6652102e-05, -1.340629e-05, -1.4925043e-06, 0.00029664068, 3.5703502e-05, -1.2303174e-05, -1.7011157e-06, 0.0002766784, 4.4005174e-05, -1.1025539e-05, -1.8807775e-06, 0.00025277736, 5.143986e-05, -9.596152e-06, -2.0288026e-06, 0.00022539719, 5.7905985e-05, -8.039967e-06, -2.1430494e-06, 0.00019504406, 6.3319065e-05, -6.383686e-06, -2.2219558e-06, 0.00016226186, 6.761283e-05, -4.655302e-06, -2.2645609e-06, 0.00012762289, 7.074005e-05, -2.8836205e-06, -2.2705158e-06, 9.171818e-05, 7.2673e-05, -1.0977758e-06, -2.2400866e-06, 5.5147735e-05, 7.340364e-05, 6.7325703e-07, -2.1741428e-06, 1.8510673e-05, 7.294342e-05, 2.4011383e-06, -2.0741388e-06, -1.7604401e-05, 7.132284e-05, 4.0586265e-06, -1.9420838e-06, -5.262873e-05, 6.8590605e-05, 5.620015e-06, -1.7805023e-06, -8.602226e-05, 6.481261e-05, 7.061542e-06, -1.5923865e-06, -0.000117281874, 6.007052e-05, 8.361757e-06, -1.3811418e-06, -0.00014594894, 5.4460226e-05, 9.501849e-06, -1.1505241e-06, -0.00017161595, 4.8090023e-05, 1.0465924e-05, -9.045725e-07, -0.00019393222, 4.1078627e-05, 1.1241232e-05, -6.475384e-07, -0.00021260865, 3.3553064e-05, 1.1818332e-05, -3.8381037e-07, -0.00022742117, 2.5646408e-05, 1.2191206e-05, -1.1783818e-07, -0.0002382134, 1.7495518e-05, 1.23573145e-05, 1.4594347e-07, -0.00024489776, 9.238686e-06, 1.2317581e-05, 4.0319043e-07, -0.00024745576, 1.0133339e-06, 1.2076334e-05, 6.497219e-07, -0.00024593686, -7.046252e-06, 1.1641178e-05, 8.815902e-07, -0.00024045652, -1.481109e-05, 1.1022821e-05, 1.0951446e-06, -0.00023119285, -2.215956e-05, 1.0234844e-05, 1.287091e-06, -0.00021838261, -2.8979288e-05, 9.293433e-06, 1.4545428e-06, -0.00020231603, -3.516886e-05, 8.217064e-06, 1.5950659e-06, -0.00018333098, -4.0639312e-05, 7.0261517e-06, 1.7067146e-06, -0.00016180646, -4.5315388e-05, 5.7426832e-06, 1.7880577e-06, -0.00013815545, -4.9136554e-05, 4.389815e-06, 1.8381979e-06, -0.00011281736, -5.2057734e-05, 2.991463e-06, 1.8567788e-06, -8.625015e-05, -5.4049786e-05, 1.571888e-06, 1.8439844e-06, -5.8922342e-05, -5.5099677e-05, 1.552773e-07, 1.8005284e-06, -3.1304942e-05, -5.521042e-05, -1.234664e-06, 1.7276353e-06, -3.863511e-06, -5.440071e-05, -2.5751076e-06, 1.6270119e-06, 2.2949533e-05, -5.2704294e-05, -3.844475e-06, 1.5008111e-06, 4.8702248e-05, -5.0169147e-05, -5.022784e-06, 1.351589e-06, 7.299001e-05, -4.685635e-05, -6.091961e-06, 1.1822551e-06, 9.5441756e-05, -4.2838827e-05, -7.036117e-06, 9.960171e-07, 0.00011572555, -3.819987e-05, -7.841781e-06, 7.96321e-07, 0.00013355333, -3.3031523e-05, -8.498087e-06, 5.8678893e-07, 0.00014868495, -2.7432841e-05, -8.996914e-06, 3.7115348e-07, 0.00016093111, -2.1508078e-05, -9.332981e-06, 1.5319195e-07, 0.00017015559, -1.5364798e-05, -9.503879e-06, -6.333968e-08, 0.00017627634, -9.111979e-06, -9.510066e-06, -2.7477122e-07, 0.00017926583, -2.8581278e-06, -9.354809e-06, -4.775805e-07, 0.0001791502, 3.2905689e-06, -9.044071e-06, -6.684519e-07, 0.00017600782, 9.232012e-06, -8.586366e-06, -8.4433054e-07, 0.00016996665, 1.4869858e-05, -7.992561e-06, -1.0024712e-06, 0.00016120113, 2.0115047e-05, -7.2756475e-06, -1.1404807e-06, 0.0001499281, 2.4887187e-05, -6.450476e-06, -1.256354e-06, 0.00013640216, 2.9115756e-05, -5.533468e-06, -1.3485029e-06, 0.00012091052, 3.274111e-05, -4.5422994e-06, -1.4157764e-06, 0.00010376727, 3.571529e-05, -3.495574e-06, -1.4574739e-06, 8.530748e-05, 3.8002585e-05, -2.4124809e-06, -1.4733498e-06, 6.5880915e-05, 3.9579925e-05, -1.312453e-06, -1.4636101e-06, 4.5845678e-05, 4.0436986e-05, -2.1482376e-07, -1.4289019e-06, 2.5561856e-05, 4.0576113e-05, 8.615063e-07, -1.3702935e-06, 5.385265e-06, 4.0012004e-05, 1.8983899e-06, -1.28925e-06, -1.4338623e-05, 3.8771206e-05, 2.8787344e-06, -1.1875999e-06, -3.3280427e-05, 3.6891386e-05, 3.7867792e-06, -1.0674974e-06, -5.1132196e-05, 3.442045e-05, 4.6083446e-06, -9.31379e-07, -6.761229e-05, 3.1415482e-05, 5.331048e-06, -7.8191624e-07, -8.246964e-05, 2.7941562e-05, 5.944487e-06, -6.219642e-07, -9.548748e-05, 2.4070448e-05, 6.4403775e-06, -4.5450886e-07, -0.00010648627, 1.9879188e-05, 6.8126637e-06, -2.8261215e-07, -0.00011532605, 1.5448655e-05, 7.0575747e-06, -1.0935682e-07, -0.00012190792, 1.086205e-05, 7.173647e-06, 6.2207974e-08, -0.00012617487, 6.2033896e-06, 7.161705e-06, 2.2911972e-07, -0.00012811176, 1.5560229e-06, 7.0247993e-06, 3.885531e-07, -0.00012774469, -2.9988225e-06, 6.76811e-06, 5.378674e-07, -0.00012513953, -7.3834203e-06, 6.398811e-06, 6.746493e-07, -0.000120399905, -1.1524835e-05, 5.9259046e-06, 7.96752e-07, -0.00011366442, -1.5356103e-05, 5.360026e-06, 9.0232743e-07, -0.00010510346, -1.8817278e-05, 4.713222e-06, 9.898541e-07, -9.4915464e-05, -2.1856336e-05, 3.9987094e-06, 1.0581577e-06, -8.332271e-05, -2.4429924e-05, 3.2306175e-06, 1.1064254e-06, -7.0566864e-05, -2.6503923e-05, 2.42372e-06, 1.1342138e-06, -5.6904282e-05, -2.8053862e-05, 1.5931603e-06, 1.1414497e-06, -4.2601067e-05, -2.9065124e-05, 7.5417444e-07, 1.1284247e-06, -2.7928161e-05, -2.9532996e-05, -7.818002e-08, 1.0957832e-06, -1.3156416e-05, -2.9462524e-05, -8.8928823e-07, 1.0445041e-06, 1.4482314e-06, -2.8868213e-05, -1.6652284e-06, 9.758777e-07, 1.562936e-05, -2.7773556e-05, -2.3930056e-06, 8.9147625e-07, 2.9144427e-05, -2.621041e-05, -3.060763e-06, 7.9312133e-07, 4.1768744e-05, -2.4218249e-05, -3.6579706e-06, 6.828461e-07, 5.32991e-05, -2.1843282e-05, -4.1755848e-06, 5.628556e-07, 6.3556865e-05, -1.9137478e-05, -4.6061787e-06, 4.3548374e-07, 7.239062e-05, -1.6157512e-05, -4.944042e-06, 3.0314965e-07, 7.9678226e-05, -1.296364e-05, -5.1852458e-06, 1.6831255e-07, 8.532833e-05, -9.618542e-06, -5.3276785e-06, 3.342723e-08, 8.928128e-05, -6.1861397e-06, -5.371042e-06, -9.909978e-08, 9.1509464e-05, -2.730425e-06, -5.3168214e-06, -2.2695231e-07, 9.201702e-05, 6.8569426e-07, -5.168221e-06, -3.4794425e-07, 9.0839065e-05, 4.0014997e-06, -4.9300693e-06, -4.6005619e-07, 8.804029e-05, 7.1595086e-06, -4.6087002e-06, -5.6146837e-07, 8.371312e-05, 1.0106435e-05, -4.2118054e-06, -6.5058947e-07, 7.7975405e-05, 1.2794058e-05, -3.7482685e-06, -7.2608077e-07, 7.096766e-05, 1.51799795e-05, -3.2279802e-06, -7.86875e-07, 6.285003e-05, 1.7228254e-05, -2.661638e-06, -8.3219066e-07, 5.3798878e-05, 1.8909906e-05, -2.0605369e-06, -8.6154023e-07, 4.4003267e-05, 2.0203282e-05, -1.4363524e-06, -8.747332e-07, 3.3661185e-05, 2.109429e-05, -8.009219e-07, -8.718737e-07, 2.297576e-05, 2.1576489e-05, -1.6602695e-07, -8.533529e-07, 1.2151434e-05, 2.1651016e-05, 4.5681873e-07, -8.1983643e-07, 1.3902205e-06, 2.1326414e-05, 1.056572e-06, -7.722467e-07, -9.111928e-06, 2.0618303e-05, 1.6228506e-06, -7.1174145e-07, -1.916855e-05, 1.954894e-05, 2.1461078e-06, -6.396881e-07, -2.8605858e-05, 1.8146657e-05, 2.6177875e-06, -5.576349e-07, -3.726562e-05, 1.6445221e-05, 3.030459e-06, -4.6727934e-07, -4.5007695e-05, 1.448309e-05, 3.3779293e-06, -3.7043466e-07, -5.1712177e-05, 1.2302602e-05, 3.6553279e-06, -2.6899448e-07, -5.7281126e-05, 9.949122e-06, 3.859169e-06, -1.6489703e-07, -6.1639854e-05, 7.470142e-06, 3.987385e-06, -6.008913e-08, -6.473777e-05, 4.9143637e-06, 4.0393347e-06, 4.3509356e-08, -6.6548724e-05, 2.330779e-06, 4.0157865e-06, 1.440398e-07, -6.707097e-05, -2.322336e-07, 3.9188717e-06, 2.397374e-07, -6.632661e-05, -2.727783e-06, 3.7520183e-06, 3.2896136e-07, -6.436064e-05, -5.111295e-06, 3.5198623e-06, 4.102223e-07, -6.12396e-05, -7.34128e-06, 3.228136e-06, 4.8220636e-07, -5.704988e-05, -9.380026e-06, 2.8835402e-06, 5.4379564e-07, -5.189563e-05, -1.1194213e-05, 2.4936026e-06, 5.9408467e-07, -4.5896457e-05, -1.2755427e-05, 2.0665202e-06, 6.323927e-07, -3.9184866e-05, -1.4040577e-05, 1.6109971e-06, 6.5827186e-07, -3.1903503e-05, -1.5032207e-05, 1.1360726e-06, 6.715103e-07, -2.420229e-05, -1.571869e-05, 6.509493e-07, 6.7213176e-07, -1.6235488e-05, -1.6094316e-05, 1.648198e-07, 6.603903e-07, -8.158729e-06, -1.615928e-05, -3.1330168e-07, 6.3676123e-07, -1.2610064e-07, -1.591953e-05, -7.747416e-07, 6.0192775e-07, 7.71268e-06, -1.5386546e-05, -1.2113197e-06, 5.5676463e-07, 1.5214951e-05, -1.4577009e-05, -1.6154895e-06, 5.0231824e-07, 2.2247606e-05, -1.3512368e-05, -1.9804643e-06, 4.3978403e-07, 2.868936e-05, -1.2218351e-05, -2.3003258e-06, 3.7048167e-07, 3.4432735e-05, -1.07243895e-05, -2.5701174e-06, 2.9582839e-07, 3.9385777e-05, -9.062992e-06, -2.7859137e-06, 2.1731096e-07, 4.347341e-05, -7.2690787e-06, -2.9448724e-06, 1.3645717e-07, 4.6638488e-05, -5.3792764e-06, -3.0452657e-06, 5.4806844e-08, 4.8842445e-05, -3.431205e-06, -3.0864876e-06, -2.6116663e-08, 5.0065628e-05, -1.4627515e-06, -3.0690437e-06, -1.0483414e-07, 5.0307255e-05, 4.886368e-07, -2.994518e-06, -1.799369e-07, 4.9585e-05, 2.3866428e-06, -2.8655218e-06, -2.5011127e-07, 4.793429e-05, 4.1967323e-06, -2.6856248e-06, -3.1416099e-07, 4.540724e-05, 5.88676e-06, -2.4592691e-06, -3.7102683e-07, 4.2071322e-05, 7.4275194e-06, -2.191669e-06, -4.1980354e-07, 3.8007787e-05, 8.793228e-06, -1.8886984e-06, -4.597535e-07, 3.3309818e-05, 9.961934e-06, -1.556769e-06, -4.9031695e-07, 2.8080553e-05, 1.091585e-05, -1.2026999e-06, -5.11119e-07, 2.2430933e-05, 1.1641598e-05, -8.3358253e-07, -5.219729e-07, 1.6477446e-05, 1.21303665e-05, -4.5664385e-07, -5.228796e-07, 1.0339824e-05, 1.23779855e-05, -7.9108844e-08, -5.1402446e-07, 4.138731e-06, 1.2384904e-05, 2.9193384e-07, -4.9576994e-07, -2.0065343e-06, 1.215609e-05, 6.496611e-07, -4.6864557e-07, -7.98025e-06, 1.1700845e-05, 9.87637e-07, -4.333348e-07, -1.3672376e-05, 1.1032538e-05, 1.2999253e-06, -3.906596e-07, -1.8980505e-05, 1.0168278e-05, 1.5811897e-06, -3.415623e-07, -2.3811644e-05, 9.128512e-06, 1.8267821e-06, -2.8708595e-07, -2.808376e-05, 7.936575e-06, 2.0328146e-06, -2.2835302e-07, -3.1727115e-05, 6.618195e-06, 2.1962185e-06, -1.6654303e-07, -3.4685316e-05, 5.2009636e-06, 2.314784e-06, -1.0286963e-07, -3.6916124e-05, 3.713776e-06, 2.3871862e-06, -3.8557374e-08, -3.8391958e-05, 2.1862647e-06, 2.4129906e-06, 2.5181173e-08, -3.9100112e-05, 6.4822814e-07, 2.3926455e-06, 8.716774e-08, -3.9042712e-05, -8.70934e-07, 2.3274554e-06, 1.4627956e-07, -3.823636e-05, -2.342765e-06, 2.2195406e-06, 2.0146919e-07, -3.6711557e-05, -3.7402674e-06, 2.0717814e-06, 2.517825e-07, -3.4511824e-05, -5.038384e-06, 1.8877496e-06, 2.9637468e-07, -3.1692645e-05, -6.214431e-06, 1.6716281e-06, 3.3452383e-07, -2.8320166e-05, -7.248476e-06, 1.4281212e-06, 3.6564208e-07, -2.4469746e-05, -8.123664e-06, 1.1623565e-06, 3.89284e-07, -2.0224345e-05, -8.826472e-06, 8.7978043e-07, 4.0515212e-07, -1.567281e-05, -9.346904e-06, 5.8605065e-07, 4.1309983e-07, -1.09080775e-05, -9.678604e-06, 2.8692546e-07, 4.1313106e-07, -6.0253424e-06, -9.818912e-06, -1.1845466e-08, 4.053976e-07, -1.1202042e-06, -9.768842e-06, -3.0462908e-07, 3.901933e-07, 3.7131454e-06, -9.532992e-06, -5.8601216e-07, 3.6794606e-07, 8.38368e-06, -9.11939e-06, -8.508988e-07, 3.392073e-07, 1.2805202e-05, -8.539277e-06, -1.0945998e-06, 3.0463937e-07, 1.6897882e-05, -7.806834e-06, -1.3129135e-06, 2.6500112e-07, 2.0589652e-05, -6.938863e-06, -1.5021946e-06, 2.2113198e-07, 2.3817425e-05, -5.9544136e-06, -1.659413e-06, 1.7393484e-07, 2.6528118e-05, -4.8743877e-06, -1.7821992e-06, 1.243579e-07, 2.8679478e-05, -3.7211096e-06, -1.8688759e-06, 7.337623e-08, 3.0240672e-05, -2.5178747e-06, -1.918477e-06, 2.1973078e-08, 3.1192667e-05, -1.2884959e-06, -1.9307531e-06, -2.8878702e-08, 3.1528372e-05, -5.6842556e-08, -1.9061621e-06, -7.8234585e-08, 3.1252544e-05, 1.1536112e-06, -1.8458483e-06, -1.2519553e-07, 3.03815e-05, 2.3202217e-06, -1.7516077e-06, -1.6892389e-07, 2.894257e-05, 3.4215889e-06, -1.6258431e-06, -2.0865801e-07, 2.6973406e-05, 4.437937e-06, -1.4715074e-06, -2.4372503e-07, 2.4521065e-05, 5.3514605e-06, -1.2920383e-06, -2.735519e-07, 2.164095e-05, 6.1466203e-06, -1.0912846e-06, -2.9767418e-07, 1.8395613e-05, 6.810402e-06, -8.7342687e-07, -3.1574282e-07, 1.4853441e-05, 7.332512e-06, -6.428926e-07, -3.275287e-07, 1.10872525e-05, 7.705526e-06, -4.0426863e-07, -3.3292451e-07, 7.172846e-06, 7.924974e-06, -1.6221205e-07, -3.3194476e-07, 3.1875018e-06, 7.989379e-06, 7.863867e-08, -3.247233e-07, -7.915006e-07, 7.900224e-06, 3.1375046e-07, -3.115085e-07, -4.688351e-06, 7.661875e-06, 5.387791e-07, -2.9265678e-07, -8.430117e-06, 7.2814523e-06, 7.496474e-07, -2.6862392e-07, -1.1948078e-05, 6.7686383e-06, 9.426174e-07, -2.3995463e-07, -1.5178949e-05, 6.135456e-06, 1.1143544e-06, -2.0727096e-07, -1.8065988e-05, 5.396e-06, 1.2619826e-06, -1.7125919e-07, -2.0559957e-05, 4.5661336e-06, 1.3831312e-06, -1.3265583e-07, -2.2619923e-05, 3.6631589e-06, 1.4759702e-06, -9.223296e-08, -2.4213892e-05, 2.705464e-06, 1.5392351e-06, -5.078315e-08, -2.5319265e-05, 1.7121589e-06, 1.572241e-06, -9.104239e-09, -2.5923093e-05, 7.0270056e-07, 1.5748852e-06, 3.2015688e-08, -2.6022171e-05, -3.0347928e-07, 1.5476394e-06, 7.181289e-08, -2.5622929e-05, -1.287341e-06, 1.4915302e-06, 1.0956186e-07, -2.4741137e-05, -2.2305894e-06, 1.4081108e-06, 1.4458821e-07, -2.3401466e-05, -3.116007e-06, 1.2994226e-06, 1.762805e-07, -2.163686e-05, -3.9277597e-06, 1.167948e-06, 2.0410044e-07, -1.9487774e-05, -4.6516734e-06, 1.0165566e-06, 2.2759187e-07, -1.7001285e-05, -5.2754713e-06, 8.4844424e-07, 2.4638777e-07, -1.4230091e-05, -5.788976e-06, 6.670677e-07, 2.6021561e-07, -1.1231426e-05, -6.1842643e-06, 4.7607486e-07, 2.6890086e-07, -8.065888e-06, -6.4557794e-06, 2.7923318e-07, 2.723685e-07, -4.7962562e-06, -6.6003963e-06, 8.035655e-08, 2.7064283e-07, -1.486253e-06, -6.6174393e-06, -1.1676697e-07, 2.6384507e-07, 1.8006667e-06, -6.5086547e-06, -3.084461e-07, 2.5218972e-07, 5.0025137e-06, -6.2781373e-06, -4.911539e-07, 2.359787e-07, 8.05991e-06, -5.9322147e-06, -6.615916e-07, 2.1559434e-07, 1.0917169e-05, -5.4792886e-06, -8.167464e-07, 1.9149074e-07, 1.3523284e-05, -4.9296464e-06, -9.539435e-07, 1.6418414e-07, 1.5832818e-05, -4.295232e-06, -1.0708909e-06, 1.3424207e-07, 1.7806671e-05, -3.5893959e-06, -1.1657154e-06, 1.0227193e-07, 1.941271e-05, -2.8266206e-06, -1.2369916e-06, 6.890892e-08, 2.0626268e-05, -2.0222278e-06, -1.2837605e-06, 3.480361e-08, 2.143049e-05, -1.1920772e-06, -1.3055406e-06, 6.0956007e-10, 2.1816513e-05, -3.5225867e-07, -1.3023282e-06, -3.3029014e-08, 2.1783524e-05, 4.812144e-07, -1.2745897e-06, -6.548915e-08, 2.1338628e-05, 1.2927053e-06, -1.2232455e-06, -9.618044e-08, 2.0496598e-05, 2.0672421e-06, -1.1496448e-06, -1.2455557e-07, 1.9279467e-05, 2.790789e-06, -1.0555334e-06, -1.501198e-07, 1.7716e-05, 3.450495e-06, -9.430141e-07, -1.7243944e-07, 1.584105e-05, 4.0349164e-06, -8.145016e-07, -1.9114883e-07, 1.369479e-05, 4.5342103e-06, -6.726722e-07, -2.0595614e-07, 1.1321889e-05, 4.940292e-06, -5.204086e-07, -2.1664762e-07, 8.7705885e-06, 5.2469613e-06, -3.6074326e-07, -2.230902e-07, 6.091738e-06, 5.449987e-06, -1.9679844e-07, -2.2523274e-07, 3.337804e-06, 5.5471555e-06, -3.1726362e-08, -2.2310557e-07, 5.6184854e-07, 5.5382793e-06, 1.3135045e-07, -2.1681858e-07, -2.1834733e-06, 5.42517e-06, 2.893973e-07, -2.0655787e-07, -4.8468987e-06, 5.21157e-06, 4.395228e-07, -1.9258094e-07, -7.3795e-06, 4.9030546e-06, 5.7903077e-07, -1.7521076e-07, -9.735567e-06, 4.5068937e-06, 7.054677e-07, -1.5482858e-07, -1.1873417e-05, 4.031892e-06, 8.166647e-07, -1.3186587e-07, -1.3756115e-05, 3.488198e-06, 9.1077374e-07, -1.0679541e-07, -1.535209e-05, 2.8870916e-06, 9.862971e-07, -8.012172e-08, -1.6635651e-05, 2.2407557e-06, 1.0421095e-06, -5.2371135e-08, -1.7587372e-05, 1.5620321e-06, 1.0774737e-06, -2.4081587e-08, -1.8194361e-05, 8.641707e-07, 1.0920477e-06, 4.2076684e-09, -1.8450402e-05, 1.6057416e-07, 1.0858846e-06, 3.1966152e-08, -1.8355964e-05, -5.3545574e-07, 1.059426e-06, 5.8681955e-08, -1.791809e-05, -1.2109659e-06, 1.0134868e-06, 8.3871015e-08, -1.7150163e-05, -1.8535899e-06, 9.492341e-07, 1.07085704e-07, -1.607156e-05, -2.4517694e-06, 8.6816004e-07, 1.2792263e-07, -1.4707189e-05, -2.9949601e-06, 7.7204817e-07, 1.4602945e-07, -1.3086937e-05, -3.4738111e-06, 6.629357e-07, 1.6111065e-07, -1.1245037e-05, -3.880323e-06, 5.430712e-07, 1.7293212e-07, -9.219358e-06, -4.2079773e-06, 4.1486925e-07, 1.8132452e-07, -7.0506335e-06, -4.4518324e-06, 2.808623e-07, 1.8618549e-07, -4.7816607e-06, -4.6085947e-06, 1.4365173e-07, 1.8748035e-07, -2.4564627e-06, -4.676652e-06, 5.8578706e-09, 1.8524176e-07, -1.1944607e-07, -4.65608e-06, -1.2992929e-07, 1.7956795e-07, 2.1854369e-06, -4.5486117e-06, -2.6119807e-07, 1.7061983e-07, 4.4155036e-06, -4.357581e-06, -3.8556084e-07, 1.5861703e-07, 6.530122e-06, -4.0878344e-06, -5.0079683e-07, 1.4383275e-07, 8.491439e-06, -3.745618e-06, -6.048907e-07, 1.2658786e-07, 1.0265044e-05, -3.3384367e-06, -6.960675e-07, 1.07244134e-07, 1.1820564e-05, -2.8748964e-06, -7.728215e-07, 8.619676e-08};
endpackage
`endif
