`ifndef data/Coefficients_FIR12_SV_
`define data/Coefficients_FIR12_SV_
package data/Coefficients_FIR12;
	localparam N = 4;
	localparam OSR = 12;
	localparam real hf[0:1999] = {0.00013426498, -4.9124017e-05, 1.7975931e-06, 7.7123175e-08, 0.00010967693, -4.915521e-05, 2.252349e-06, 5.4354526e-08, 8.518222e-05, -4.8751986e-05, 2.6926682e-06, 2.7658853e-08, 6.0995677e-05, -4.7924703e-05, 3.113002e-06, -2.5885363e-09, 3.7325797e-05, -4.668822e-05, 3.5081152e-06, -3.596963e-08, 1.437256e-05, -4.5061675e-05, 3.8731423e-06, -7.2029614e-08, -7.674623e-06, -4.3068212e-05, 4.20364e-06, -1.1028309e-07, -2.8638853e-05, -4.073464e-05, 4.495633e-06, -1.5022056e-07, -4.835748e-05, -3.8091097e-05, 4.7456556e-06, -1.9131505e-07, -6.6683664e-05, -3.5170637e-05, 4.950782e-06, -2.3302891e-07, -8.348776e-05, -3.2008826e-05, 5.108656e-06, -2.7482048e-07, -9.86584e-05, -2.8643286e-05, 5.2175074e-06, -3.1615085e-07, -0.00011210349, -2.5113257e-05, 5.276167e-06, -3.5649023e-07, -0.00012375083, -2.145911e-05, 5.284069e-06, -3.9532458e-07, -0.00013354862, -1.7721877e-05, 5.241251e-06, -4.3216122e-07, -0.0001414656, -1.3942781e-05, 5.1483435e-06, -4.6653489e-07, -0.00014749111, -1.0162762e-05, 5.0065532e-06, -4.980127e-07, -0.00015163478, -6.42202e-06, 4.817643e-06, -5.261991e-07, -0.00015392606, -2.759572e-06, 4.583901e-06, -5.507401e-07, -0.00015441353, 7.871683e-07, 4.308108e-06, -5.713269e-07, -0.00015316399, 4.1827884e-06, 3.993496e-06, -5.876991e-07, -0.00015026134, 7.3942438e-06, 3.6437077e-06, -5.996472e-07, -0.0001458054, 1.0391191e-05, 3.2627433e-06, -6.070144e-07, -0.0001399104, 1.3146283e-05, 2.854914e-06, -6.0969785e-07, -0.0001327034, 1.5635434e-05, 2.4247845e-06, -6.076492e-07, -0.00012432267, 1.7838025e-05, 1.9771173e-06, -6.0087456e-07, -0.00011491592, 1.9737088e-05, 1.5168157e-06, -5.8943357e-07, -0.000104638355, 2.1319423e-05, 1.0488639e-06, -5.7343834e-07, -9.365084e-05, 2.257569e-05, 5.7826946e-07, -5.5305145e-07, -8.211792e-05, 2.3500439e-05, 1.1000523e-07, -5.2848327e-07, -7.020592e-05, 2.4092109e-05, -3.5104782e-07, -4.999891e-07, -5.808097e-05, 2.4352963e-05, -8.001546e-07, -4.6786565e-07, -4.5907123e-05, 2.4289007e-05, -1.2327786e-06, -4.3244722e-07, -3.384453e-05, 2.390984e-05, -1.6446301e-06, -3.9410114e-07, -2.2047687e-05, 2.322849e-05, -2.0317125e-06, -3.532234e-07, -1.066375e-05, 2.2261183e-05, -2.3903626e-06, -3.1023364e-07, 1.689847e-07, 2.1027123e-05, -2.7172882e-06, -2.6557012e-07, 1.0322505e-05, 1.954819e-05, -3.0095994e-06, -2.1968441e-07, 1.968035e-05, 1.7848655e-05, -3.2648356e-06, -1.730362e-07, 2.8138724e-05, 1.5954853e-05, -3.4809868e-06, -1.2608793e-07, 3.560744e-05, 1.3894836e-05, -3.65651e-06, -7.9299475e-08, 4.2010703e-05, 1.1698021e-05, -3.7903378e-06, -3.312308e-08, 4.7287678e-05, 9.394823e-06, -3.881885e-06, 1.20016965e-08, 5.139292e-05, 7.016283e-06, -3.931046e-06, 5.565275e-08, 5.4296575e-05, 4.5937004e-06, -3.93819e-06, 9.7429925e-08, 5.5984437e-05, 2.1582607e-06, -3.904146e-06, 1.3695919e-07, 5.645778e-05, -2.59322e-07, -3.830189e-06, 1.7389642e-07, 5.5733046e-05, -2.6291552e-06, -3.7180175e-06, 2.0793094e-07, 5.3841355e-05, -4.9225e-06, -3.5697249e-06, 2.3878832e-07, 5.0827828e-05, -7.1120844e-06, -3.3877711e-06, 2.6623303e-07, 4.675081e-05, -9.172396e-06, -3.1749487e-06, 2.9007043e-07, 4.16809e-05, -1.1079947e-05, -2.9343437e-06, 3.1014832e-07, 3.569988e-05, -1.28135125e-05, -2.6692965e-06, 3.263579e-07, 2.8899538e-05, -1.4354335e-05, -2.3833597e-06, 3.3863438e-07, 2.1380387e-05, -1.5686304e-05, -2.0802527e-06, 3.4695688e-07, 1.3250306e-05, -1.6796095e-05, -1.7638173e-06, 3.513481e-07, 4.623113e-06, -1.7673276e-05, -1.4379715e-06, 3.5187307e-07, -4.3828954e-06, -1.8310377e-05, -1.1066631e-06, 3.486379e-07, -1.3646438e-05, -1.870293e-05, -7.7382435e-07, 3.4178785e-07, -2.3044748e-05, -1.8849465e-05, -4.4332685e-07, 3.315049e-07, -3.2455067e-05, -1.8751478e-05, -1.1893848e-07, 3.1800516e-07, -4.1756113e-05, -1.8413355e-05, 1.9571803e-07, 3.0153583e-07, -5.0829505e-05, -1.7842283e-05, 4.9720404e-07, 2.823717e-07, -5.9561116e-05, -1.704811e-05, 7.823013e-07, 2.6081173e-07, -6.784239e-05, -1.6043183e-05, 1.048045e-06, 2.3717516e-07, -7.5571515e-05, -1.4842162e-05, 1.291753e-06, 2.1179738e-07, -8.265456e-05, -1.34618185e-05, 1.5110523e-06, 1.8502608e-07, -8.900645e-05, -1.1920787e-05, 1.7039002e-06, 1.5721683e-07, -9.455183e-05, -1.0239331e-05, 1.8686025e-06, 1.2872903e-07, -9.922587e-05, -8.439066e-06, 2.0038258e-06, 9.992165e-08, -0.00010297478, -6.542694e-06, 2.1086075e-06, 7.114919e-08, -0.000105756364, -4.573715e-06, 2.1823598e-06, 4.27577e-08, -0.000107540305, -2.5561385e-06, 2.2248694e-06, 1.5080946e-08, -0.000108308355, -5.141956e-07, 2.236294e-06, -1.1563163e-08, -0.00010805439, 1.5279481e-06, 2.217153e-06, -3.6875946e-08, -0.00010678427, 3.5464745e-06, 2.1683152e-06, -6.0581e-08, -0.000104515646, 5.5181854e-06, 2.090983e-06, -8.242701e-08, -0.00010127755, 7.4207633e-06, 1.9866714e-06, -1.0219011e-07, -9.7109885e-05, 9.233017e-06, 1.8571858e-06, -1.19676e-07, -9.2062844e-05, 1.0935116e-05, 1.7045952e-06, -1.3472165e-07, -8.619614e-05, 1.250879e-05, 1.5312035e-06, -1.4719652e-07, -7.957819e-05, 1.3937526e-05, 1.3395185e-06, -1.5700354e-07, -7.2285184e-05, 1.520673e-05, 1.1322194e-06, -1.6407958e-07, -6.440013e-05, 1.6303866e-05, 9.1212195e-07, -1.6839554e-07, -5.6011726e-05, 1.7218566e-05, 6.821435e-07, -1.6995605e-07, -4.721333e-05, 1.7942724e-05, 4.452671e-07, -1.687988e-07, -3.8101745e-05, 1.8470546e-05, 2.0450557e-07, -1.6499347e-07, -2.8776105e-05, 1.879859e-05, -3.71344e-08, -1.586403e-07, -1.933667e-05, 1.8925755e-05, -2.766871e-07, -1.4986844e-07, -9.883665e-06, 1.8853274e-05, -5.112619e-07, -1.3883376e-07, -5.161338e-07, 1.858465e-05, -7.380757e-07, -1.2571665e-07, 8.669189e-06, 1.812558e-05, -9.544837e-07, -1.1071944e-07, 1.7578946e-05, 1.7483864e-05, -1.1580076e-06, -9.406355e-08, 2.6124177e-05, 1.6669272e-05, -1.3463628e-06, -7.598662e-08, 3.422127e-05, 1.5693402e-05, -1.5174804e-06, -5.673939e-08, 4.179284e-05, 1.4569521e-05, -1.669529e-06, -3.658251e-08, 4.876851e-05, 1.331238e-05, -1.8009314e-06, -1.578331e-08, 5.508561e-05, 1.1938023e-05, -1.910379e-06, 5.3874767e-09, 6.0689777e-05, 1.0463577e-05, -1.9968431e-06, 2.6658975e-08, 6.553543e-05, 8.907045e-06, -2.0595814e-06, 4.776336e-08, 6.9586175e-05, 7.2870757e-06, -2.0981424e-06, 6.843896e-08, 7.281505e-05, 5.6227427e-06, -2.1123658e-06, 8.843324e-08, 7.520467e-05, 3.9333177e-06, -2.1023802e-06, 1.0750564e-07, 7.6747325e-05, 2.2380445e-06, -2.068596e-06, 1.2543022e-07, 7.744484e-05, 5.559175e-07, -2.0116956e-06, 1.4199803e-07, 7.730846e-05, -1.0945329e-06, -1.932623e-06, 1.5701937e-07, 7.635852e-05, -2.695445e-06, -1.8325662e-06, 1.7032569e-07, 7.462406e-05, -4.2298216e-06, -1.7129411e-06, 1.8177117e-07, 7.21424e-05, -5.6817107e-06, -1.5753701e-06, 1.9123415e-07, 6.895852e-05, -7.036372e-06, -1.4216607e-06, 1.9861817e-07, 6.512443e-05, -8.280426e-06, -1.2537811e-06, 2.0385264e-07, 6.069849e-05, -9.401988e-06, -1.0738347e-06, 2.068933e-07, 5.5744564e-05, -1.0390773e-05, -8.840334e-07, 2.0772241e-07, 5.0331266e-05, -1.1238196e-05, -6.866704e-07, 2.0634833e-07, 4.453106e-05, -1.1937436e-05, -4.840919e-07, 2.0280527e-07, 3.8419366e-05, -1.2483488e-05, -2.7866915e-07, 1.9715227e-07, 3.207364e-05, -1.2873186e-05, -7.277051e-08, 1.8947229e-07, 2.5572472e-05, -1.3105215e-05, 1.31266e-07, 1.7987074e-07, 1.8994639e-05, -1.3180086e-05, 3.311594e-07, 1.6847399e-07, 1.2418219e-05, -1.3100107e-05, 5.2471125e-07, 1.5542756e-07, 5.919696e-06, -1.286932e-05, 7.098298e-07, 1.4089409e-07, -4.268843e-07, -1.2493429e-05, 8.8455255e-07, 1.250512e-07, -6.5507234e-06, -1.1979699e-05, 1.0470668e-06, 1.0808921e-07, -1.2385025e-05, -1.1336854e-05, 1.1957283e-06, 9.020873e-08, -1.7867693e-05, -1.0574948e-05, 1.3290776e-06, 7.161814e-08, -2.294196e-05, -9.705219e-06, 1.4458537e-06, 5.253109e-08, -2.7556945e-05, -8.739949e-06, 1.5450061e-06, 3.3163914e-08, -3.1668136e-05, -7.6923e-06, 1.6257023e-06, 1.3733093e-08, -3.5237783e-05, -6.576144e-06, 1.6873352e-06, -5.547255e-09, -3.8235223e-05, -5.405895e-06, 1.7295255e-06, -2.4467816e-08, -4.0637085e-05, -4.1963294e-06, 1.7521227e-06, -4.282643e-08, -4.242745e-05, -2.9624093e-06, 1.7552034e-06, -6.04303e-08, -4.3597895e-05, -1.7191086e-06, 1.7390659e-06, -7.709811e-08, -4.4147433e-05, -4.812366e-07, 1.7042239e-06, -9.266187e-08, -4.408242e-05, 7.367289e-07, 1.6513966e-06, -1.0696872e-07, -4.3416323e-05, 1.9208044e-06, 1.581497e-06, -1.198824e-07, -4.216946e-05, 3.0576537e-06, 1.4956184e-06, -1.3128457e-07, -4.0368614e-05, 4.134731e-06, 1.3950184e-06, -1.4107589e-07, -3.8046615e-05, 5.1404136e-06, 1.2811022e-06, -1.4917686e-07, -3.5241854e-05, 6.0641187e-06, 1.1554031e-06, -1.5552841e-07, -3.1997726e-05, 6.8964105e-06, 1.0195636e-06, -1.6009227e-07, -2.8362047e-05, 7.6290876e-06, 8.7531413e-07, -1.6285102e-07, -2.4386396e-05, 8.255259e-06, 7.244514e-07, -1.6380802e-07, -2.012547e-05, 8.769397e-06, 5.688172e-07, -1.6298695e-07, -1.5636371e-05, 9.1673855e-06, 4.102756e-07, -1.6043128e-07, -1.09779085e-05, 9.446534e-06, 2.506917e-07, -1.5620341e-07, -6.2098743e-06, 9.605592e-06, 9.190987e-08, -1.5038361e-07, -1.3923286e-06, 9.644734e-06, -6.4267304e-08, -1.4306886e-07, 3.4151067e-06, 9.565535e-06, -2.1609894e-07, -1.3437136e-07, 8.153938e-06, 9.370926e-06, -3.61925e-07, -1.2441713e-07, 1.27674675e-05, 9.06514e-06, -5.0018406e-07, -1.1334416e-07, 1.7201422e-05, 8.6536365e-06, -6.294295e-07, -1.01300735e-07, 2.1404547e-05, 8.14302e-06, -7.483446e-07, -8.844353e-08, 2.5329156e-05, 7.5409416e-06, -8.557551e-07, -7.493563e-08, 2.8931634e-05, 6.8559925e-06, -9.506405e-07, -6.094457e-08, 3.2172866e-05, 6.0975885e-06, -1.0321435e-06, -4.6640334e-08, 3.5018624e-05, 5.2758464e-06, -1.0995764e-06, -3.2193338e-08, 3.7439895e-05, 4.401454e-06, -1.1524268e-06, -1.777247e-08, 3.9413117e-05, 3.4855357e-06, -1.19036e-06, -3.543172e-09, 4.0920375e-05, 2.5395161e-06, -1.2132202e-06, 1.0334412e-08, 4.194951e-05, 1.5749823e-06, -1.221029e-06, 2.3707189e-08, 4.249417e-05, 6.035457e-07, -1.2139822e-06, 3.6430755e-08, 4.255379e-05, -3.6329317e-07, -1.1924438e-06, 4.837091e-08, 4.213349e-05, -1.3142766e-06, -1.1569404e-06, 5.940504e-08, 4.1243944e-05, -2.2385163e-06, -1.1081505e-06, 6.94233e-08, 3.9901144e-05, -3.1256145e-06, -1.0468954e-06, 7.832969e-08, 3.8126134e-05, -3.9657757e-06, -9.741264e-07, 8.6042895e-08, 3.594469e-05, -4.7499107e-06, -8.909117e-07, 9.249699e-08, 3.3386932e-05, -5.4697316e-06, -7.984223e-07, 9.7641895e-08, 3.0486905e-05, -6.117833e-06, -6.9791633e-07, 1.014437e-07, 2.7282123e-05, -6.6877633e-06, -5.907229e-07, 1.0388479e-07, 2.3813078e-05, -7.1740856e-06, -4.7822556e-07, 1.0496369e-07, 2.0122709e-05, -7.5724224e-06, -3.6184537e-07, 1.0469487e-07, 1.6255875e-05, -7.879488e-06, -2.4302366e-07, 1.03108256e-07, 1.2258806e-05, -8.093112e-06, -1.2320504e-07, 1.00248606e-07, 8.178529e-06, -8.212241e-06, -3.820437e-09, 9.6174745e-08, 4.062324e-06, -8.236934e-06, 1.13729186e-07, 9.095863e-08, -4.283608e-08, -8.168347e-06, 2.280886e-07, 8.468425e-08, -4.090821e-06, -8.008697e-06, 3.3796326e-07, 7.74465e-08, -8.036867e-06, -7.761217e-06, 4.4213328e-07, 6.93498e-08, -1.183807e-05, -7.4301074e-06, 5.394664e-07, 6.050681e-08, -1.5453854e-05, -7.0204683e-06, 6.2892946e-07, 5.103687e-08, -1.8846404e-05, -6.538223e-06, 7.095989e-07, 4.1064588e-08, -2.1981054e-05, -5.9900403e-06, 7.806696e-07, 3.0718237e-08, -2.482664e-05, -5.383241e-06, 8.4146194e-07, 2.012822e-08, -2.7355805e-05, -4.725704e-06, 8.914279e-07, 9.425508e-09, -2.9545245e-05, -4.025767e-06, 9.301548e-07, -1.2598905e-09, -3.137592e-05, -3.292118e-06, 9.573683e-07, -1.1800431e-08, -3.2833203e-05, -2.5336944e-06, 9.729329e-07, -2.2072472e-08, -3.3906967e-05, -1.759571e-06, 9.768507e-07, -3.1957654e-08, -3.4591645e-05, -9.788552e-07, 9.692602e-07, -4.134418e-08, -3.48862e-05, -2.0057973e-07, 9.504314e-07, -5.0128005e-08, -3.479408e-05, 5.663997e-07, 9.2076056e-07, -5.8213924e-08, -3.432309e-05, 1.3135045e-06, 8.807639e-07, -6.5516524e-08, -3.3485238e-05, 2.0325276e-06, 8.3106903e-07, -7.196099e-08, -3.2296517e-05, 2.7157218e-06, 7.7240634e-07, -7.748384e-08, -3.077667e-05, 3.3558824e-06, 7.055983e-07, -8.2033424e-08, -2.8948893e-05, 3.9464207e-06, 6.3154863e-07, -8.557036e-08, -2.6839498e-05, 4.48143e-06, 5.5123024e-07, -8.8067765e-08, -2.4477575e-05, 4.955743e-06, 4.656731e-07, -8.951135e-08, -2.1894599e-05, 5.364978e-06, 3.759509e-07, -8.989939e-08, -1.9124036e-05, 5.705577e-06, 2.8316816e-07, -8.924251e-08, -1.6200916e-05, 5.9748345e-06, 1.8844688e-07, -8.75634e-08, -1.3161405e-05, 6.1709106e-06, 9.291303e-08, -8.489627e-08, -1.0042372e-05, 6.292841e-06, -2.3163729e-09, -8.128634e-08, -6.8809495e-06, 6.340532e-06, -9.614614e-08, -7.678906e-08, -3.7141008e-06, 6.314747e-06, -1.8751525e-07, -7.1469344e-08, -5.7819847e-07, 6.217085e-06, -2.754086e-07, -6.5400634e-08, 2.4913857e-06, 6.049943e-06, -3.5886794e-07, -5.8663908e-08, 5.4606708e-06, 5.8164806e-06, -4.3700206e-07, -5.134661e-08, 8.297437e-06, 5.520568e-06, -5.08996e-07, -4.3541533e-08, 1.0971562e-05, 5.1667275e-06, -5.741192e-07, -3.5345646e-08, 1.3455338e-05, 4.7600743e-06, -6.317326e-07, -2.6858908e-08, 1.5723748e-05, 4.3062428e-06, -6.8129435e-07, -1.8183052e-08, 1.7754708e-05, 3.8113158e-06, -7.223647e-07, -9.420371e-09, 1.9529267e-05, 3.2817456e-06, -7.546092e-07, -6.725389e-10, 2.103178e-05, 2.724273e-06, -7.778008e-07, 7.960574e-09, 2.2250024e-05, 2.1458443e-06, -7.9182087e-07, 1.6382023e-08, 2.3175287e-05, 1.5535279e-06, -7.966585e-07, 2.4498855e-08, 2.3802402e-05, 9.544302e-07, -7.9240914e-07, 3.222313e-08, 2.4129746e-05, 3.5561303e-07, -7.792713e-07, 3.947285e-08, 2.41592e-05, -2.3598747e-07, -7.575429e-07, 4.617281e-08, 2.3896067e-05, -8.1363885e-07, -7.27616e-07, 5.2255363e-08, 2.3348948e-05, -1.3708867e-06, -6.899706e-07, 5.7661047e-08, 2.2529586e-05, -1.9016246e-06, -6.4516786e-07, 6.233918e-08, 2.145268e-05, -2.400159e-06, -5.9384206e-07, 6.6248276e-08, 2.0135658e-05, -2.8612676e-06, -5.36692e-07, 6.935635e-08, 1.859843e-05, -3.280252e-06, -4.7447202e-07, 7.164119e-08, 1.6863112e-05, -3.6529834e-06, -4.079822e-07, 7.3090376e-08, 1.4953742e-05, -3.9759407e-06, -3.3805844e-07, 7.370132e-08, 1.2895951e-05, -4.2462393e-06, -2.655621e-07, 7.348111e-08, 1.0716654e-05, -4.461656e-06, -1.9136974e-07, 7.244624e-08, 8.443707e-06, -4.6206424e-06, -1.1636257e-07, 7.062232e-08, 6.1055703e-06, -4.7223302e-06, -4.141635e-08, 6.8043576e-08, 3.730968e-06, -4.766532e-06, 3.260873e-08, 6.4752335e-08, 1.3485509e-06, -4.75373e-06, 1.0487771e-07, 6.079839e-08, -1.0134366e-06, -4.6850596e-06, 1.7459004e-07, 5.623832e-08, -3.3274757e-06, -4.562284e-06, 2.4098833e-07, 5.11347e-08, -5.5670807e-06, -4.3877667e-06, 3.033663e-07, 4.5555286e-08, -7.707088e-06, -4.1644284e-06, 3.610761e-07, 3.9572154e-08, -9.723927e-06, -3.895709e-06, 4.1353488e-07, 3.326079e-08, -1.15958655e-05, -3.5855153e-06, 4.6023024e-07, 2.6699158e-08, -1.3303231e-05, -3.238169e-06, 5.0072515e-07, 1.996677e-08, -1.48286035e-05, -2.8583506e-06, 5.346617e-07, 1.314373e-08, -1.615698e-05, -2.4510373e-06, 5.617637e-07, 6.3098113e-09, -1.7275908e-05, -2.0214409e-06, 5.8183883e-07, -4.564637e-10, -1.8175586e-05, -1.5749441e-06, 5.9477907e-07, -7.0787065e-09, -1.8848932e-05, -1.1170346e-06, 6.005608e-07, -1.3483507e-08, -1.9291623e-05, -6.532397e-07, 5.992435e-07, -1.9601229e-08, -1.9502093e-05, -1.8906177e-07, 5.9096766e-07, -2.5366752e-08, -1.948151e-05, 2.700851e-07, 5.759519e-07, -3.072014e-08, -1.9233712e-05, 7.189366e-07, 5.5448896e-07, -3.560725e-08, -1.876512e-05, 1.1524363e-06, 5.2694116e-07, -3.9980257e-08, -1.8084624e-05, 1.5657911e-06, 4.9373494e-07, -4.3798096e-08, -1.7203425e-05, 1.9545223e-06, 4.5535492e-07, -4.702682e-08, -1.6134885e-05, 2.3145117e-06, 4.1233733e-07, -4.9639873e-08, -1.489432e-05, 2.6420444e-06, 3.6526276e-07, -5.1618272e-08, -1.3498795e-05, 2.9338432e-06, 3.1474897e-07, -5.2950696e-08, -1.1966899e-05, 3.1871018e-06, 2.6144284e-07, -5.3633475e-08, -1.0318504e-05, 3.3995066e-06, 2.0601249e-07, -5.3670522e-08, -8.574506e-06, 3.5692574e-06, 1.4913931e-07, -5.3073144e-08, -6.756573e-06, 3.6950785e-06, 9.150964e-08, -5.185978e-08, -4.8868797e-06, 3.7762247e-06, 3.3806906e-08, -5.005569e-08, -2.9878381e-06, 3.812482e-06, -2.329634e-08, -4.7692517e-08, -1.0818374e-06, 3.8041599e-06, -7.914597e-08, -4.4807837e-08, 8.0901765e-07, 3.7520797e-06, -1.3311355e-07, -4.1444608e-08, 2.6631562e-06, 3.6575564e-06, -1.8460318e-07, -3.7650587e-08, 4.4597846e-06, 3.5223748e-06, -2.3305786e-07, -3.3477697e-08, 6.179112e-06, 3.3487618e-06, -2.7796526e-07, -2.8981354e-08, 7.802566e-06, 3.139352e-06, -3.1886293e-07, -2.4219762e-08, 9.312984e-06, 2.8971513e-06, -3.5534273e-07, -1.9253203e-08, 1.0694792e-05, 2.6254954e-06, -3.870548e-07, -1.41432945e-08, 1.1934158e-05, 2.3280056e-06, -4.1371035e-07, -8.952257e-09, 1.301912e-05, 2.0085429e-06, -4.3508436e-07, -3.7421835e-09, 1.3939699e-05, 1.6711579e-06, -4.5101672e-07, 1.4256752e-09, 1.4687975e-05, 1.3200414e-06, -4.6141324e-07, 6.4916086e-09, 1.5258151e-05, 9.594742e-07, -4.6624558e-07, 1.139811e-08, 1.564658e-05, 5.9377464e-07, -4.655504e-07, 1.6090505e-08, 1.5851776e-05, 2.2724912e-07, -4.5942787e-07, 2.0517534e-08, 1.5874388e-05, -1.3585822e-07, -4.4803951e-07, 2.46319e-08, 1.5717165e-05, -4.9141335e-07, -4.316052e-07, 2.8390728e-08, 1.5384887e-05, -8.3543836e-07, -4.1039968e-07, 3.175601e-08, 1.488427e-05, -1.1641552e-06, -3.847484e-07, 3.469495e-08, 1.4223866e-05, -1.4740253e-06, -3.5502302e-07, 3.7180254e-08, 1.3413924e-05, -1.7617879e-06, -3.2163618e-07, 3.9190365e-08, 1.246625e-05, -2.0244916e-06, -2.850361e-07, 4.0709605e-08, 1.1394041e-05, -2.2595245e-06, -2.4570082e-07, 4.1728267e-08, 1.0211711e-05, -2.4646383e-06, -2.0413209e-07, 4.224262e-08, 8.934701e-06, -2.637968e-06, -1.6084921e-07, 4.2254854e-08, 7.579287e-06, -2.7780475e-06, -1.163827e-07, 4.1772964e-08, 6.1623746e-06, -2.8838201e-06, -7.126793e-08, 4.081054e-08, 4.7012963e-06, -2.954643e-06, -2.6038887e-08, 3.9386535e-08, 3.2136004e-06, -2.9902883e-06, 1.8777998e-08, 3.7524952e-08, 1.7168471e-06, -2.9909393e-06, 6.2669855e-08, 3.5254473e-08, 2.2840403e-07, -2.9571802e-06, 1.05143066e-07, 3.2608053e-08, -1.2347514e-06, -2.8899838e-06, 1.4572868e-07, 2.9622475e-08, -2.656221e-06, -2.790693e-06, 1.839874e-07, 2.6337844e-08, -4.020367e-06, -2.6609994e-06, 2.1951423e-07, 2.2797076e-08, -5.3124786e-06, -2.5029176e-06, 2.5194257e-07, 1.9045359e-08, -6.518927e-06, -2.3187565e-06, 2.809478e-07, 1.512958e-08, -7.6273054e-06, -2.111088e-06, 3.0625037e-07, 1.1097757e-08, -8.626552e-06, -1.8827121e-06, 3.276183e-07, 6.9984707e-09, -9.507054e-06, -1.6366218e-06, 3.44869e-07, 2.8802822e-09, -1.0260735e-05, -1.3759638e-06, 3.5787062e-07, -1.2088235e-09, -1.0881122e-05, -1.1040007e-06, 3.6654274e-07, -5.2219864e-09, -1.1363397e-05, -8.2407036e-07, 3.7085647e-07, -9.113995e-09, -1.17044165e-05, -5.3954653e-07, 3.7083376e-07, -1.2841783e-08, -1.1902729e-05, -2.537991e-07, 3.665465e-07, -1.6364893e-08, -1.19585575e-05, 2.984493e-08, 3.5811473e-07, -1.9645904e-08, -1.1873768e-05, 3.0813928e-07, 3.4570454e-07, -2.2650813e-08, -1.1651824e-05, 5.7795455e-07, 3.2952522e-07, -2.5349369e-08, -1.1297717e-05, 8.3631244e-07, 3.0982628e-07, -2.7715366e-08, -1.0817882e-05, 1.0804179e-06, 2.8689377e-07, -2.972688e-08, -1.0220101e-05, 1.3076881e-06, 2.6104647e-07, -3.136645e-08, -9.513387e-06, 1.5157791e-06, 2.3263149e-07, -3.262121e-08, -8.707863e-06, 1.7026088e-06, 2.0201998e-07, -3.3482948e-08, -7.814621e-06, 1.8663766e-06, 1.6960222e-07, -3.394815e-08, -6.845581e-06, 2.0055795e-06, 1.3578291e-07, -3.4017937e-08, -5.813336e-06, 2.1190249e-06, 1.0097623e-07, -3.369799e-08, -4.7309973e-06, 2.2058382e-06, 6.5600815e-08, -3.2998404e-08, -3.6120318e-06, 2.2654688e-06, 3.0074894e-08, -3.19335e-08, -2.470101e-06, 2.2976901e-06, -5.1885602e-09, -3.0521583e-08, -1.3188992e-06, 2.3025973e-06, -3.9786546e-08, -2.8784674e-08, -1.7199385e-07, 2.2806e-06, -7.333052e-08, -2.6748188e-08, 9.573292e-07, 2.2324134e-06, -1.0545065e-07, -2.4440578e-08, 2.056215e-06, 2.1590433e-06, -1.3579982e-07, -2.1892962e-08, 3.112381e-06, 2.0617713e-06, -1.6405721e-07, -1.9138719e-08, 4.1142503e-06, 1.9421338e-06, -1.8993164e-07, -1.6213058e-08, 5.0510735e-06, 1.8019003e-06, -2.131644e-07, -1.31525875e-08, 5.913039e-06, 1.6430498e-06, -2.3353171e-07, -9.994863e-09, 6.6913713e-06, 1.467743e-06, -2.5084674e-07, -6.777935e-09, 7.378416e-06, 1.2782954e-06, -2.6496116e-07, -3.5399075e-09, 7.9677075e-06, 1.0771467e-06, -2.7576613e-07, -3.184874e-10, 8.454026e-06, 8.668317e-07, -2.8319306e-07, 2.8494411e-09, 8.833436e-06, 6.4994805e-07, -2.872136e-07, 5.9282312e-09, 9.10331e-06, 4.2912583e-07, -2.8783927e-07, 8.883866e-09, 9.262337e-06, 2.0699648e-07, -2.851208e-07, 1.16843255e-08, 9.3105145e-06, -1.3838067e-08, -2.7914672e-07, 1.4299923e-08, 9.249132e-06, -2.3083474e-07, -2.700418e-07, 1.6703611e-08, 9.080723e-06, -4.41538e-07, -2.5796498e-07, 1.8871251e-08, 8.809027e-06, -6.4360677e-07, -2.4310694e-07, 2.0781846e-08, 8.4389185e-06, -8.348396e-07, -2.2568727e-07, 2.2417723e-08, 7.97633e-06, -1.013198e-06, -2.0595165e-07, 2.3764692e-08, 7.428173e-06, -1.176827e-06, -1.8416834e-07, 2.481215e-08, 6.8022323e-06, -1.3240742e-06, -1.6062482e-07, 2.5553138e-08, 6.1070673e-06, -1.4535045e-06, -1.3562409e-07, 2.5984367e-08, 5.351898e-06, -1.5639142e-06, -1.094809e-07, 2.610619e-08, 4.546485e-06, -1.6543402e-06, -8.2517914e-08, 2.5922537e-08, 3.7010093e-06, -1.7240675e-06, -5.5061825e-08, 2.5440816e-08, 2.825947e-06, -1.7726331e-06, -2.74395e-08, 2.4671758e-08, 1.9319414e-06, -1.7998278e-06, 2.5803368e-11, 2.3629244e-08, 1.0296783e-06, -1.805693e-06, 2.7018132e-08, 2.233009e-08, 1.2976001e-07, -1.7905174e-06, 5.323237e-08, 2.0793799e-08, -7.5741497e-07, -1.7548286e-06, 7.83776e-08, 1.9042291e-08, -1.6217699e-06, -1.6993832e-06, 1.0218024e-07, 1.7099612e-08, -2.4536614e-06, -1.6251545e-06, 1.243869e-07, 1.4991617e-08, -3.243983e-06, -1.5333167e-06, 1.44767e-07, 1.2745634e-08, -3.9842625e-06, -1.4252289e-06, 1.6311506e-07, 1.03901305e-08, -4.6667506e-06, -1.3024157e-06, 1.7925264e-07, 7.954359e-09, -5.2844953e-06, -1.1665467e-06, 1.9302996e-07, 5.4680056e-09, -5.8314126e-06, -1.0194148e-06, 2.0432718e-07, 2.960839e-09, -6.3023413e-06, -8.629132e-07, 2.1305522e-07, 4.623623e-10, -6.6930857e-06, -6.990124e-07, 2.1915633e-07, -1.998524e-09, -7.0004508e-06, -5.297349e-07, 2.2260423e-07, -4.393847e-09, -7.2222597e-06, -3.5713194e-07, 2.234038e-07, -6.696871e-09, -7.3573647e-06, -1.8325862e-07, 2.2159064e-07, -8.882386e-09, -7.40564e-06, -1.01502735e-08, 2.1722998e-07, -1.0926977e-08, -7.3679694e-06, 1.6020091e-07, 2.1041555e-07, -1.280926e-08, -7.2462153e-06, 3.258682e-07, 2.0126794e-07, -1.4510102e-08, -7.0431843e-06, 4.850115e-07, 1.8993275e-07, -1.6012798e-08, -6.7625765e-06, 6.358975e-07, 1.7657851e-07, -1.7303236e-08, -6.408928e-06, 7.7691743e-07, 1.6139433e-07, -1.8369999e-08, -5.9875456e-06, 9.066042e-07, 1.445873e-07, -1.920447e-08, -5.50443e-06, 1.0236466e-06, 1.263799e-07, -1.9800869e-08, -4.9661962e-06, 1.1269021e-06, 1.07007054e-07, -2.0156282e-08, -4.3799864e-06, 1.215407e-06, 8.671322e-08, -2.0270647e-08, -3.7533775e-06, 1.288385e-06, 6.574943e-08, -2.01467e-08, -3.0942876e-06, 1.3452525e-06, 4.437024e-08, -1.9789896e-08, -2.4108767e-06, 1.3856223e-06, 2.28307e-08, -1.9208306e-08, -1.7114489e-06, 1.4093055e-06, 1.3834331e-09, -1.8412473e-08, -1.0043543e-06, 1.4163087e-06, -1.972429e-08, -1.7415251e-08, -2.9789044e-07, 1.4068324e-06, -4.0253312e-08, -1.6231615e-08, 3.9979207e-07, 1.3812643e-06, -5.997523e-08, -1.4878451e-08, 1.080782e-06, 1.3401719e-06, -7.867485e-08, -1.3374327e-08, 1.7374947e-06, 1.2842931e-06, -9.615249e-08, -1.1739254e-08, 2.362755e-06, 1.2145244e-06, -1.12226e-07, -9.99442e-09, 2.9498726e-06, 1.1319082e-06, -1.2673257e-07, -8.161933e-09, 3.492712e-06, 1.0376182e-06, -1.3953034e-07, -6.264544e-09, 3.985754e-06, 9.329429e-07, -1.5049966e-07, -4.325372e-09, 4.4241497e-06, 8.1927e-07, -1.5954407e-07, -2.3676316e-09, 4.8037637e-06, 6.9806754e-07, -1.6659106e-07, -4.1435996e-10, 5.121212e-06, 5.7086595e-07, -1.7159255e-07, 1.5118462e-09, 5.373887e-06, 4.3923941e-07, -1.745249e-07, 3.3890863e-09, 5.559975e-06, 3.0478648e-07, -1.7538893e-07, 5.196398e-09, 5.6784647e-06, 1.6911157e-07, -1.7420939e-07, 6.913984e-09, 5.7291436e-06, 3.380595e-08, -1.710343e-07, 8.523424e-09, 5.712588e-06, -9.957028e-08, -1.6593397e-07, 1.000786e-08, 5.6301433e-06, -2.2950583e-07, -1.5899988e-07, 1.1352173e-08, 5.4838933e-06, -3.5455486e-07, -1.5034318e-07, 1.2543124e-08, 5.2766272e-06, -4.733526e-07, -1.4009314e-07, 1.35694735e-08, 5.011792e-06, -5.846299e-07, -1.2839526e-07, 1.4422085e-08, 4.6934424e-06, -6.872262e-07, -1.1540938e-07, 1.5093987e-08, 4.326185e-06, -7.8010106e-07, -1.0130757e-07, 1.5580424e-08, 3.9151128e-06, -8.623445e-07, -8.627191e-08, 1.587887e-08, 3.4657407e-06, -9.3318494e-07, -7.049221e-08, 1.5989023e-08, 2.9839332e-06, -9.91996e-07, -5.4163714e-08, 1.5912766e-08, 2.4758301e-06, -1.0383012e-06, -3.7484686e-08, 1.5654114e-08, 1.9477716e-06, -1.0717773e-06, -2.0654124e-08, 1.5219124e-08, 1.4062213e-06, -1.0922547e-06, -3.8694035e-09, 1.4615798e-08, 8.5768846e-07, -1.0997175e-06, 1.2675972e-08, 1.3853953e-08, 3.086531e-07, -1.0943008e-06, 2.8794547e-08, 1.2945072e-08, -2.3450959e-07, -1.0762866e-06, 4.430698e-08, 1.1902151e-08, -7.6560093e-07, -1.046098e-06, 5.904399e-08, 1.07395195e-08, -1.2786675e-06, -1.0042918e-06, 7.284814e-08, 9.472648e-09, -1.7680661e-06, -9.515502e-07, 8.5575465e-08, 8.117954e-09, -2.2285237e-06, -8.886704e-07, 9.709691e-08, 6.6925936e-09, -2.6551927e-06, -8.165533e-07, 1.0729957e-07, 5.2142486e-09, -3.0436986e-06, -7.3619185e-07, 1.1608772e-07, 3.7009165e-09, -3.3901845e-06, -6.4865736e-07, 1.2338364e-07, 2.1706932e-09, -3.6913455e-06, -5.550862e-07, 1.2912822e-07, 6.415631e-10, -3.944458e-06, -4.5666536e-07, 1.3328129e-07, -8.688073e-10, -4.1474023e-06, -3.546179e-07, 1.3582181e-07, -2.3432691e-09, -4.298675e-06, -2.5018807e-07, 1.3674774e-07, -3.765381e-09, -4.397398e-06, -1.4462663e-07, 1.3607581e-07, -5.119587e-09, -4.443317e-06, -3.9176268e-08, 1.3384093e-07, -6.3913816e-09, -4.436793e-06, 6.4942704e-08, 1.3009554e-07, -7.567461e-09, -4.3787904e-06, 1.665461e-07, 1.2490865e-07, -8.635855e-09, -4.2708525e-06, 2.6449896e-07, 1.1836482e-07, -9.586044e-09, -4.1150765e-06, 3.5772788e-07, 1.1056285e-07, -1.0409056e-08, -3.9140773e-06, 4.452323e-07, 1.0161446e-07, -1.1097543e-08, -3.6709498e-06, 5.26095e-07, 9.164274e-08, -1.1645841e-08, -3.3892256e-06, 5.994913e-07, 8.0780524e-08, -1.2050004e-08, -3.0728231e-06, 6.646967e-07, 6.9168706e-08, -1.230782e-08, -2.7259969e-06, 7.210943e-07, 5.695448e-08, -1.2418811e-08, -2.3532814e-06, 7.681793e-07, 4.42895e-08, -1.2384206e-08, -1.959435e-06, 8.0556356e-07, 3.1328064e-08, -1.2206895e-08, -1.5493806e-06, 8.329778e-07, 1.8225295e-08, -1.1891376e-08, -1.1281453e-06, 8.5027267e-07, 5.135308e-09, -1.1443665e-08, -7.0080125e-07, 8.574188e-07, -7.790542e-09, -1.0871206e-08, -2.724054e-07, 8.545047e-07, -2.040537e-08, -1.0182761e-08, 1.5205823e-07, 8.41734e-07, -3.2568387e-08, -9.388285e-09, 5.6773547e-07, 8.19421e-07, -4.414642e-08, -8.498788e-09, 9.699559e-07, 7.879853e-07, -5.5015335e-08, -7.526194e-09, 1.3542835e-06, 7.479449e-07, -6.506131e-08, -6.483184e-09, 1.716565e-06, 6.999089e-07, -7.4181976e-08, -5.383038e-09, 2.0529717e-06, 6.4456856e-07, -8.228743e-08, -4.2394706e-09, 2.36004e-06, 5.826882e-07, -8.930103e-08, -3.0664649e-09, 2.6347043e-06, 5.1509477e-07, -9.516009e-08, -1.8781057e-09, 2.8743257e-06, 4.4266764e-07, -9.981635e-08, -6.8841594e-10, 3.0767164e-06, 3.6632716e-07, -1.0323628e-07, 4.8880555e-10, 3.2401558e-06, 2.8702343e-07, -1.05401256e-07, 1.6401397e-09, 3.3634042e-06, 2.0572494e-07, -1.06307475e-07, 2.7526954e-09, 3.4457078e-06, 1.2340685e-07, -1.05965796e-07, 3.8142507e-09, 3.4868e-06, 4.1039677e-08, -1.0440132e-07, 4.8133812e-09, 3.4868958e-06, -4.0421888e-08, -1.01652894e-07, 5.739581e-09, 3.4466816e-06, -1.2004975e-07, -9.7772414e-08, 6.583366e-09, 3.3672984e-06, -1.969527e-07, -9.282399e-08, 7.3363675e-09, 3.250322e-06, -2.7028614e-07, -8.688303e-08, 7.991411e-09, 3.0977371e-06, -3.3926105e-07, -8.003514e-08, 8.542577e-09, 2.9119071e-06, -4.0315217e-07, -7.2374995e-08, 8.985249e-09, 2.6955406e-06, -4.6130543e-07, -6.400504e-08, 9.316144e-09, 2.4516537e-06, -5.131441e-07, -5.5034256e-08, 9.53333e-09, 2.183531e-06, -5.5817435e-07, -4.5576684e-08, 9.6362225e-09, 1.8946821e-06, -5.9598955e-07, -3.57501e-08, 9.6255715e-09, 1.5887973e-06, -6.262734e-07, -2.5674563e-08, 9.503425e-09, 1.2697021e-06, -6.4880214e-07, -1.5470972e-08, 9.27309e-09, 9.413105e-07, -6.634457e-07, -5.2596714e-09, 8.939068e-09, 6.0757816e-07, -6.701672e-07, 4.8409365e-09, 8.506984e-09, 2.7245602e-07, -6.6902237e-07, 1.47157335e-08, 7.983502e-09, -6.015555e-08, -6.6015696e-07, 2.425416e-08, 7.3762334e-09, -3.864509e-07, -6.438037e-07, 3.3351416e-08, 6.6936265e-09, -7.0276155e-07, -6.2027794e-07, 4.190958e-08, 5.944862e-09, -1.0055966e-06, -5.8997296e-07, 4.9838622e-08, 5.1397278e-09, -1.2916796e-06, -5.533537e-07, 5.7057317e-08, 4.2885e-09, -1.5579836e-06, -5.109505e-07, 6.3494035e-08, 3.401815e-09, -1.8017615e-06, -4.6335154e-07, 6.90874e-08, 2.4905382e-09, -2.020573e-06, -4.1119546e-07, 7.3786836e-08, 1.5656364e-09, -2.2123081e-06, -3.5516274e-07, 7.755298e-08, 6.380493e-10, -2.375206e-06, -2.959673e-07, 8.035793e-08, -2.8143765e-10, -2.5078689e-06, -2.3434765e-07, 8.2185366e-08, -1.1823145e-09, -2.6092728e-06, -1.710579e-07, 8.3030585e-08, -2.054464e-09, -2.678773e-06, -1.06858806e-07, 8.290033e-08, -2.8882718e-09, -2.7161043e-06, -4.25088e-08, 8.1812495e-08, -3.67473e-09, -2.7213791e-06, 2.1244709e-08, 7.979579e-08, -4.4055297e-09, -2.6950786e-06, 8.367381e-08, 7.688919e-08, -5.073146e-09, -2.6380412e-06, 1.440782e-07, 7.314129e-08, -5.670912e-09, -2.5514473e-06, 2.017928e-07, 6.860964e-08, -6.193082e-09, -2.4367994e-06, 2.561949e-07, 6.335987e-08, -6.6348798e-09, -2.2958993e-06, 3.0671066e-07, 5.7464828e-08, -6.992541e-09, -2.1308224e-06, 3.5282082e-07, 5.1003614e-08, -7.2633384e-09, -1.943889e-06, 3.9406595e-07, 4.4060535e-08, -7.4455935e-09, -1.7376329e-06, 4.3005068e-07, 3.6724067e-08, -7.538683e-09, -1.5147697e-06, 4.6044713e-07, 2.908575e-08, -7.543022e-09, -1.2781605e-06, 4.849977e-07, 2.1239083e-08, -7.460051e-09, -1.0307779e-06, 5.035169e-07, 1.32784e-08, -7.292191e-09, -7.7566847e-07, 5.15892e-07, 5.2977662e-09, -7.0428072e-09, -5.1591746e-07, 5.220835e-07, -2.6100968e-09, -6.716151e-09, -2.546114e-07, 5.2212397e-07, -1.0354873e-08, -6.317297e-09, 5.1971494e-09, 5.161168e-07, -1.7849652e-08, -5.8520677e-09, 2.605245e-07, 5.042337e-07, -2.5011877e-08, -5.3269584e-09};
	localparam real hb[0:1999] = {0.00015872756, -4.865276e-05, 1.3341992e-06, 9.5637695e-08, 0.00018284425, -4.774062e-05, 8.6815066e-07, 1.0962415e-07, 0.0002063954, -4.6391695e-05, 4.0554585e-07, 1.1886612e-07, 0.00022916467, -4.4615e-05, -4.7474618e-08, 1.2320822e-07, 0.00025094146, -4.2424464e-05, -4.848008e-07, 1.225591e-07, 0.00027152334, -3.9838804e-05, -9.00428e-07, 1.16893595e-07, 0.0002907184, -3.6881396e-05, -1.2885312e-06, 1.062542e-07, 0.00030834752, -3.358006e-05, -1.6435382e-06, 9.075168e-08, 0.00032424656, -2.9966797e-05, -1.9602016e-06, 7.05649e-08, 0.0003382684, -2.607747e-05, -2.2336678e-06, 4.5939647e-08, 0.00035028474, -2.195144e-05, -2.4595413e-06, 1.718668e-08, 0.00036018764, -1.763115e-05, -2.6339465e-06, -1.5321136e-08, 0.00036789116, -1.31616725e-05, -2.753583e-06, -5.1152586e-08, 0.00037333247, -8.590218e-06, -2.8157738e-06, -8.9822684e-08, 0.0003764727, -3.9656056e-06, -2.8185093e-06, -1.3079804e-07, 0.0003772977, 6.6228574e-07, -2.7604815e-06, -1.7350303e-07, 0.00037581843, 5.24309e-06, -2.6411105e-06, -2.1732647e-07, 0.000372071, 9.7265365e-06, -2.4605638e-06, -2.6162922e-07, 0.00036611652, 1.4063045e-05, -2.219765e-06, -3.05752e-07, 0.00035804062, 1.8204311e-05, -1.920395e-06, -3.4902368e-07, 0.00034795262, 2.2103895e-05, -1.5648823e-06, -3.9077008e-07, 0.00033598446, 2.571779e-05, -1.1563842e-06, -4.3032293e-07, 0.0003222894, 2.9004965e-05, -6.987602e-07, -4.6702863e-07, 0.0003070403, 3.192788e-05, -1.965338e-07, -5.0025744e-07, 0.00029042785, 3.445298e-05, 3.4515222e-07, -5.294122e-07, 0.0002726585, 3.655112e-05, 9.2059065e-07, -5.539371e-07, 0.00025395196, 3.8197966e-05, 1.5235717e-06, -5.7332574e-07, 0.00023453892, 3.9374336e-05, 2.147452e-06, -5.871286e-07, 0.0002146583, 4.0066472e-05, 2.7852313e-06, -5.9496074e-07, 0.00019455445, 4.026626e-05, 3.4296327e-06, -5.9650745e-07, 0.0001744744, 3.9971383e-05, 4.0731893e-06, -5.9153024e-07, 0.0001546648, 3.9185412e-05, 4.708333e-06, -5.798714e-07, 0.00013536912, 3.7917795e-05, 5.3274894e-06, -5.614574e-07, 0.00011682458, 3.618383e-05, 5.9231675e-06, -5.3630146e-07, 9.925935e-05, 3.4004497e-05, 6.4880574e-06, -5.0450507e-07, 8.288971e-05, 3.1406293e-05, 7.0151214e-06, -4.6625803e-07, 6.791738e-05, 2.8420927e-05, 7.497684e-06, -4.218376e-07, 5.4527005e-05, 2.5084999e-05, 7.929522e-06, -3.7160615e-07, 4.2883756e-05, 2.1439593e-05, 8.304945e-06, -3.1600783e-07, 3.313126e-05, 1.7529814e-05, 8.618875e-06, -2.5556398e-07, 2.538969e-05, 1.3404268e-05, 8.866912e-06, -1.9086733e-07, 1.9754154e-05, 9.114508e-06, 9.045406e-06, -1.2257519e-07, 1.6293374e-05, 4.714413e-06, 9.151499e-06, -5.140169e-08, 1.5048682e-05, 2.5955836e-07, 9.183181e-06, 2.1890996e-08, 1.603334e-05, -4.1934586e-06, 9.139315e-06, 9.6502184e-08, 1.9232195e-05, -8.587703e-06, 9.019665e-06, 1.7160292e-07, 2.460169e-05, -1.2866601e-05, 8.82491e-06, 2.4634667e-07, 3.2070217e-05, -1.6974638e-05, 8.556639e-06, 3.1988057e-07, 4.1538817e-05, -2.0858053e-05, 8.217344e-06, 3.9135682e-07, 5.288223e-05, -2.4465513e-05, 7.810396e-06, 4.5994415e-07, 6.595028e-05, -2.7748758e-05, 7.340009e-06, 5.2483927e-07, 8.056954e-05, -3.0663232e-05, 6.8111976e-06, 5.852782e-07, 9.654537e-05, -3.3168646e-05, 6.2297186e-06, 6.405467e-07, 0.00011366417, -3.522952e-05, 5.602002e-06, 6.8999105e-07, 0.00013169588, -3.681564e-05, 4.9350797e-06, 7.330269e-07, 0.00015039672, -3.7902468e-05, 4.2364977e-06, 7.6914864e-07, 0.0001695122, -3.8471495e-05, 3.5142255e-06, 7.979363e-07, 0.00018878006, -3.8510498e-05, 2.7765573e-06, 8.1906256e-07, 0.0002079336, -3.8013724e-05, 2.03201e-06, 8.322979e-07, 0.00022670485, -3.698201e-05, 1.2892147e-06, 8.375145e-07, 0.00024482794, -3.5422814e-05, 5.5680937e-07, 8.346887e-07, 0.00026204233, -3.335013e-05, -1.5667254e-07, 8.239023e-07, 0.00027809615, -3.0784387e-05, -8.429109e-07, 8.05342e-07, 0.00029274923, -2.7752207e-05, -1.4939062e-06, 7.792975e-07, 0.00030577628, -2.4286099e-05, -2.1020835e-06, 7.4615843e-07, 0.00031696958, -2.0424097e-05, -2.6603911e-06, 7.06409e-07, 0.0003261418, -1.620931e-05, -3.162393e-06, 6.6062245e-07, 0.00033312826, -1.1689395e-05, -3.602354e-06, 6.0945285e-07, 0.00033778916, -6.916003e-06, -3.9753154e-06, 5.536269e-07, 0.00034001138, -1.9441345e-06, -4.277161e-06, 4.939339e-07, 0.00033970998, 3.1685208e-06, -4.5046745e-06, 4.3121494e-07, 0.00033682946, 8.362296e-06, -4.6555797e-06, 3.6635137e-07, 0.0003313444, 1.3576281e-05, -4.7285757e-06, 3.0025262e-07, 0.0003232601, 1.8749075e-05, -4.7233525e-06, 2.3384334e-07, 0.00031261242, 2.381955e-05, -4.640599e-06, 1.6805059e-07, 0.00029946762, 2.8727603e-05, -4.4819935e-06, 1.0379065e-07, 0.00028392157, 3.3414915e-05, -4.250185e-06, 4.195609e-08, 0.0002660987, 3.7825674e-05, -3.948758e-06, -1.6596921e-08, 0.00024615065, 4.1907257e-05, -3.5821874e-06, -7.1060846e-08, 0.00022425433, 4.5610912e-05, -3.1557793e-06, -1.2068831e-07, 0.00020060995, 4.8892347e-05, -2.6756031e-06, -1.6480286e-07, 0.0001754387, 5.1712283e-05, -2.148412e-06, -2.0280861e-07, 0.00014898, 5.4036955e-05, -1.5815533e-06, -2.3419892e-07, 0.000121488716, 5.5838518e-05, -9.828734e-07, -2.5856366e-07, 9.323204e-05, 5.709539e-05, -3.606136e-07, -2.7559506e-07, 6.448637e-05, 5.779252e-05, 2.7669782e-07, -2.8509234e-07, 3.5533947e-05, 5.792157e-05, 9.2035805e-07, -2.8696442e-07, 6.659485e-06, 5.7481007e-05, 1.5616042e-06, -2.8123134e-07, -2.1853248e-05, 5.6476107e-05, 2.1917285e-06, -2.6802397e-07, -4.9724804e-05, 5.4918877e-05, 2.8021927e-06, -2.4758205e-07, -7.668339e-05, 5.2827898e-05, 3.3847393e-06, -2.2025071e-07, -0.0001024681, 5.022807e-05, 3.931501e-06, -1.8647545e-07, -0.00012683198, 4.7150286e-05, 4.435101e-06, -1.4679563e-07, -0.00014954495, 4.3631037e-05, 4.8887514e-06, -1.0183663e-07, -0.0001703965, 3.9711922e-05, 5.2863375e-06, -5.2300773e-08, -0.00018919804, 3.5439138e-05, 5.6225e-06, 1.0429668e-09, -0.00020578512, 3.086286e-05, 5.8926994e-06, 5.737008e-08, -0.00022001927, 2.6036625e-05, 6.0932744e-06, 1.1581253e-07, -0.00023178944, 2.101664e-05, 6.2214867e-06, 1.7547133e-07, -0.00024101326, 1.5861067e-05, 6.275553e-06, 2.354296e-07, -0.00024763774, 1.0629304e-05, 6.254664e-06, 2.9476575e-07, -0.00025163972, 5.3812287e-06, 6.1589917e-06, 3.525669e-07, -0.00025302602, 1.7646191e-07, 5.9896793e-06, 4.0794197e-07, -0.000251833, -4.926374e-06, 5.748825e-06, 4.6003439e-07, -0.00024812593, -9.870375e-06, 5.4394472e-06, 5.0803453e-07, -0.00024199794, -1.4601047e-05, 5.06544e-06, 5.511911e-07, -0.00023356875, -1.9066967e-05, 4.631516e-06, 5.8882193e-07, -0.00022298278, -2.322039e-05, 4.143141e-06, 6.2032336e-07, -0.0002104074, -2.7017819e-05, 3.6064553e-06, 6.451791e-07, -0.00019603045, -3.04205e-05, 3.0281908e-06, 6.6296684e-07, -0.00018005798, -3.3394866e-05, 2.415577e-06, 6.733644e-07, -0.00016271134, -3.5912908e-05, 1.776242e-06, 6.7615395e-07, -0.00014422451, -3.7952457e-05, 1.1181111e-06, 6.712245e-07, -0.00012484101, -3.9497412e-05, 4.4929916e-07, 6.585734e-07, -0.0001048109, -4.0537874e-05, -2.2199683e-07, 6.383058e-07, -8.4387575e-05, -4.1070194e-05, -8.8760595e-07, 6.1063264e-07, -6.382472e-05, -4.1096966e-05, -1.5394902e-06, 5.758674e-07, -4.3373195e-05, -4.0626903e-05, -2.1698486e-06, 5.3442096e-07, -2.3277991e-05, -3.9674673e-05, -2.7712174e-06, 4.8679544e-07, -3.775331e-06, -3.8260638e-05, -3.3365636e-06, 4.3357673e-07, 1.4910092e-05, -3.6410518e-05, -3.8593744e-06, 3.754255e-07, 3.2567714e-05, -3.4155015e-05, -4.333736e-06, 3.1306766e-07, 4.9003473e-05, -3.1529362e-05, -4.7544036e-06, 2.4728388e-07, 6.404195e-05, -2.8572813e-05, -5.1168663e-06, 1.7889803e-07, 7.7528246e-05, -2.5328101e-05, -5.4173947e-06, 1.0876556e-07, 8.932958e-05, -2.1840855e-05, -5.653081e-06, 3.7761243e-08, 9.933658e-05, -1.8158978e-05, -5.82187e-06, -3.3233157e-08, 0.00010746427, -1.4332024e-05, -5.9225736e-06, -1.0334121e-07, 0.00011365272, -1.04105375e-05, -5.954875e-06, -1.7170397e-07, 0.00011786738, -6.4454093e-06, -5.9193253e-06, -2.3749176e-07, 0.0001200991, -2.4872284e-06, -5.817322e-06, -2.9991543e-07, 0.00012036383, 1.4143535e-06, -5.651081e-06, -3.582368e-07, 0.00011870198, 5.211232e-06, -5.423598e-06, -4.1177861e-07, 0.00011517749, 8.857433e-06, -5.138596e-06, -4.5993295e-07, 0.000109876644, 1.2309665e-05, -4.800469e-06, -5.0216914e-07, 0.000102906604, 1.5527814e-05, -4.414215e-06, -5.380402e-07, 9.43937e-05, 1.8475406e-05, -3.9853617e-06, -5.6718784e-07, 8.448148e-05, 2.1120008e-05, -3.5198873e-06, -5.8934654e-07, 7.332865e-05, 2.3433568e-05, -3.024135e-06, -6.043461e-07, 6.110679e-05, 2.5392696e-05, -2.5047261e-06, -6.121125e-07, 4.7997935e-05, 2.6978882e-05, -1.9684699e-06, -6.1266803e-07, 3.4192155e-05, 2.8178645e-05, -1.4222705e-06, -6.061293e-07, 1.9884963e-05, 2.8983619e-05, -8.730384e-07, -5.9270457e-07, 5.2747746e-06, 2.9390565e-05, -3.2759874e-07, -5.7268966e-07, -9.439641e-06, 2.9401319e-05, 2.073946e-07, -5.464622e-07, -2.4061686e-05, 2.9022684e-05, 7.255425e-07, -5.144758e-07, -3.8399365e-05, 2.8266242e-05, 1.2207789e-06, -4.77252e-07, -5.2267627e-05, 2.7148137e-05, 1.687443e-06, -4.3537258e-07, -6.549057e-05, 2.5688767e-05, 2.1203455e-06, -3.8947033e-07, -7.790348e-05, 2.3912462e-05, 2.514826e-06, -3.4021963e-07, -8.935473e-05, 2.1847087e-05, 2.8668046e-06, -2.8832642e-07, -9.970742e-05, 1.9523637e-05, 3.172822e-06, -2.3451813e-07, -0.0001088408, 1.6975777e-05, 3.4300729e-06, -1.7953315e-07, -0.00011665157, 1.4239361e-05, 3.6364283e-06, -1.2411071e-07, -0.0001230548, 1.1351946e-05, 3.7904506e-06, -6.8980654e-08, -0.00012798459, 8.352278e-06, 3.891397e-06, -1.4853671e-08, -0.00013139469, 5.2797786e-06, 3.939214e-06, 3.7588073e-08, -0.00013325858, 2.1740386e-06, 3.9345255e-06, 8.769966e-08, -0.00013356947, -9.2568706e-07, 3.8786084e-06, 1.348815e-07, -0.00013234004, -3.980967e-06, 3.7733635e-06, 1.785866e-07, -0.00012960186, -6.9546595e-06, 3.621275e-06, 2.183269e-07, -0.00012540464, -9.811351e-06, 3.4253683e-06, 2.5367868e-07, -0.00011981532, -1.2517772e-05, 3.1891564e-06, 2.8428704e-07, -0.00011291682, -1.5043158e-05, 2.9165853e-06, 3.0986902e-07, -0.000104806786, -1.7359594e-05, 2.6119721e-06, 3.3021607e-07, -9.5596006e-05, -1.9442296e-05, 2.2799418e-06, 3.4519508e-07, -8.540686e-05, -2.1269858e-05, 1.9253594e-06, 3.5474838e-07, -7.437152e-05, -2.2824444e-05, 1.5532623e-06, 3.5889286e-07, -6.263016e-05, -2.4091938e-05, 1.1687919e-06, 3.5771788e-07, -5.032908e-05, -2.5062032e-05, 7.77124e-07, 3.5138225e-07, -3.7618734e-05, -2.5728274e-05, 3.8340252e-07, 3.4011043e-07, -2.4651872e-05, -2.6088062e-05, -7.3262543e-09, 3.2418768e-07, -1.1581571e-05, -2.61426e-05, -3.9017564e-07, 3.0395475e-07, 1.4406131e-06, -2.5896776e-05, -7.6047706e-07, 2.7980164e-07, 1.4266469e-05, -2.5359039e-05, -1.1138343e-06, 2.521611e-07, 2.675286e-05, -2.454121e-05, -1.4461725e-06, 2.215015e-07, 3.8763355e-05, -2.345825e-05, -1.7537823e-06, 1.8831948e-07, 5.0169736e-05, -2.212801e-05, -2.0333566e-06, 1.5313243e-07, 6.085338e-05, -2.0570948e-05, -2.2820234e-06, 1.1647084e-07, 7.0706476e-05, -1.880981e-05, -2.4973701e-06, 7.887061e-08, 7.9633086e-05, -1.6869304e-05, -2.6774615e-06, 4.086569e-08, 8.755005e-05, -1.4775753e-05, -2.8208524e-06, 2.9807488e-09, 9.4387695e-05, -1.2556725e-05, -2.9265918e-06, -3.427567e-08, 0.00010009037, -1.0240682e-05, -2.9942225e-06, -7.041763e-08, 0.0001046168, -7.856605e-06, -3.0237723e-06, -1.0498777e-07, 0.00010794026, -5.433634e-06, -3.0157407e-06, -1.3756268e-07, 0.000110048546, -3.000708e-06, -2.9710795e-06, -1.6775766e-07, 0.00011094382, -5.862235e-07, -2.8911684e-06, -1.9523077e-07, 0.00011064223, 1.782292e-06, -2.7777855e-06, -2.1968616e-07, 0.000109173394, 4.0784917e-06, -2.633074e-06, -2.4087666e-07, 0.00010657977, 6.277494e-06, -2.4595047e-06, -2.5860567e-07, 0.000102915816, 8.356144e-06, -2.259837e-06, -2.727281e-07, 9.824709e-05, 1.0293244e-05, -2.0370744e-06, -2.8315085e-07, 9.264923e-05, 1.2069758e-05, -1.794423e-06, -2.8983231e-07, 8.6206805e-05, 1.36689805e-05, -1.5352438e-06, -2.927812e-07, 7.901212e-05, 1.5076678e-05, -1.2630078e-06, -2.9205492e-07, 7.116396e-05, 1.6281187e-05, -9.812507e-07, -2.8775702e-07, 6.2766296e-05, 1.7273487e-05, -6.9352683e-07, -2.8003447e-07, 5.392692e-05, 1.8047243e-05, -4.0336622e-07, -2.69074e-07, 4.475613e-05, 1.8598805e-05, -1.1423196e-07, -2.5509843e-07, 3.536538e-05, 1.8927174e-05, 1.705193e-07, -2.3836239e-07, 2.5865978e-05, 1.9033956e-05, 4.4767467e-07, -2.191478e-07, 1.6367781e-05, 1.8923263e-05, 7.141992e-07, -1.9775923e-07, 6.978001e-06, 1.860161e-05, 9.672665e-07, -1.7451909e-07, -2.199989e-06, 1.8077764e-05, 1.2042864e-06, -1.4976267e-07, -1.1067724e-05, 1.736259e-05, 1.4229277e-06, -1.2383335e-07, -1.953266e-05, 1.6468866e-05, 1.621138e-06, -9.7077766e-08, -2.7509079e-05, 1.5411088e-05, 1.7971596e-06, -6.9841235e-08, -3.49189e-05, 1.4205255e-05, 1.9495396e-06, -4.246325e-08, -4.169237e-05, 1.2868649e-05, 2.0771388e-06, -1.5273379e-08, -4.776864e-05, 1.1419599e-05, 2.1791332e-06, 1.1412633e-08, -5.3096253e-05, 9.877248e-06, 2.255015e-06, 3.7296346e-08, -5.7633468e-05, 8.261315e-06, 2.3045877e-06, 6.2099765e-08, -6.1348495e-05, 6.591852e-06, 2.3279583e-06, 8.5568054e-08, -6.4219625e-05, 4.8890142e-06, 2.325527e-06, 1.0747179e-07, -6.623517e-05, 3.1728284e-06, 2.2979718e-06, 1.2760886e-07, -6.73934e-05, 1.4629718e-06, 2.2462334e-06, 1.458058e-07, -6.770229e-05, -2.2143733e-07, 2.1714952e-06, 1.6191879e-07, -6.717919e-05, -1.8620384e-06, 2.0751627e-06, 1.7583415e-07, -6.58504e-05, -3.441412e-06, 1.9588404e-06, 1.8746842e-07, -6.375067e-05, -4.943248e-06, 1.8243073e-06, 1.9676813e-07, -6.092257e-05, -6.3524963e-06, 1.6734924e-06, 2.0370904e-07, -5.741588e-05, -7.655499e-06, 1.5084481e-06, 2.0829516e-07, -5.3286825e-05, -8.840106e-06, 1.331324e-06, 2.105574e-07, -4.8597307e-05, -9.895765e-06, 1.1443404e-06, 2.1055197e-07, -4.3414086e-05, -1.08136e-05, 9.497624e-07, 2.0835857e-07, -3.780794e-05, -1.1586462e-05, 7.4987366e-07, 2.0407823e-07, -3.1852767e-05, -1.2208961e-05, 5.4695175e-07, 1.9783124e-07, -2.5624733e-05, -1.2677488e-05, 3.432443e-07, 1.8975473e-07, -1.9201354e-05, -1.2990196e-05, 1.4094579e-07, 1.8000033e-07, -1.2660636e-05, -1.3146991e-05, -5.7823364e-08, 1.6873166e-07, -6.0802004e-06, -1.3149479e-05, -2.5103694e-07, 1.5612196e-07, 4.635453e-07, -1.3000914e-05, -4.367809e-07, 1.4235155e-07, 6.896217e-06, -1.27061185e-05, -6.1326983e-07, 1.276056e-07, 1.3146218e-05, -1.2271399e-05, -7.7886136e-07, 1.1207178e-07, 1.9145455e-05, -1.1704446e-05, -9.320686e-07, 9.5938056e-08, 2.483e-05, -1.1014211e-05, -1.071571e-06, 7.939073e-08, 3.014069e-05, -1.0210796e-05, -1.1962222e-06, 6.261252e-08, 3.502368e-05, -9.30531e-06, -1.3050577e-06, 4.578083e-08, 3.943089e-05, -8.309739e-06, -1.3972984e-06, 2.9066195e-08, 4.3320437e-05, -7.236793e-06, -1.4723538e-06, 1.26309265e-08, 4.665693e-05, -6.0997604e-06, -1.5298226e-06, -3.3720955e-09, 4.941174e-05, -4.91236e-06, -1.5694919e-06, -1.8800428e-08, 5.1563176e-05, -3.6885833e-06, -1.5913345e-06, -3.35229e-08, 5.3096577e-05, -2.4425465e-06, -1.5955039e-06, -4.7420265e-08, 5.4004337e-05, -1.1883395e-06, -1.5823296e-06, -6.0385716e-08, 5.428586e-05, 6.011901e-08, -1.5523083e-06, -7.23252e-08, 5.3947442e-05, 1.2892245e-06, -1.5060965e-06, -8.315763e-08, 5.300207e-05, 2.4858207e-06, -1.4445001e-06, -9.281495e-08, 5.1469164e-05, 3.6373287e-06, -1.3684634e-06, -1.0124207e-07, 4.937427e-05, 4.7318663e-06, -1.2790574e-06, -1.08396726e-07, 4.6748683e-05, 5.7583597e-06, -1.177467e-06, -1.14249204e-07, 4.3629e-05, 6.7066435e-06, -1.0649773e-06, -1.1878201e-07, 4.005666e-05, 7.5675525e-06, -9.4295973e-07, -1.219895e-07, 3.6077425e-05, 8.332999e-06, -8.1285776e-07, -1.2387743e-07, 3.17408e-05, 8.9960395e-06, -6.761714e-07, -1.2446239e-07, 2.7099486e-05, 9.550929e-06, -5.344423e-07, -1.2377136e-07, 2.2208726e-05, 9.993164e-06, -3.8923855e-07, -1.2184111e-07, 1.7125712e-05, 1.0319511e-05, -2.421394e-07, -1.1871761e-07, 1.1908932e-05, 1.0528019e-05, -9.471996e-08, -1.1445547e-07, 6.6175194e-06, 1.0618026e-05, 5.146373e-08, -1.09117295e-07, 1.3106252e-06, 1.0590146e-05, 1.9488924e-07, -1.0277313e-07, -3.9532233e-06, 1.044625e-05, 3.3408196e-07, -9.5499765e-08, -9.116739e-06, 1.0189422e-05, 4.6762872e-07, -8.738017e-08, -1.4124476e-05, 9.8239225e-06, 5.941908e-07, -7.8502836e-08, -1.8923394e-05, 9.355123e-06, 7.12516e-07, -6.896113e-08, -2.3463408e-05, 8.7894405e-06, 8.2145004e-07, -5.8852645e-08, -2.769788e-05, 8.134254e-06, 9.1994724e-07, -4.8278533e-08, -3.158409e-05, 7.3978226e-06, 1.0070794e-06, -3.734283e-08, -3.508365e-05, 6.589184e-06, 1.0820445e-06, -2.6151731e-08, -3.816285e-05, 5.7180537e-06, 1.1441736e-06, -1.4812911e-08, -4.0792995e-05, 4.7947137e-06, 1.1929363e-06, -3.434746e-09, -4.295065e-05, 3.8299004e-06, 1.2279463e-06, 7.874425e-09, -4.4617835e-05, 2.8346828e-06, 1.2489633e-06, 1.9007091e-08, -4.578216e-05, 1.8203448e-06, 1.2558955e-06, 2.985737e-08, -4.6436908e-05, 7.982599e-07, 1.2487999e-06, 4.0321837e-08, -4.658104e-05, -2.2022978e-07, 1.2278805e-06, 5.030033e-08, -4.6219167e-05, -1.2239361e-06, 1.1934867e-06, 5.969683e-08, -4.536142e-05, -2.2019437e-06, 1.1461084e-06, 6.8420285e-08, -4.4023294e-05, -3.1437269e-06, 1.0863711e-06, 7.638545e-08, -4.2225434e-05, -4.0392583e-06, 1.0150286e-06, 8.3513704e-08, -3.999335e-05, -4.879118e-06, 9.3295534e-07, 8.973389e-08, -3.735708e-05, -5.6545873e-06, 8.411367e-07, 9.4983065e-08, -3.4350847e-05, -6.3577427e-06, 7.4065804e-07, 9.920721e-08, -3.1012598e-05, -6.981534e-06, 6.326937e-07, 1.02361966e-07, -2.7383587e-05, -7.519858e-06, 5.1849366e-07, 1.04413154e-07, -2.350786e-05, -7.967619e-06, 3.9937026e-07, 1.0533739e-07, -1.9431758e-05, -8.320775e-06, 2.7668403e-07, 1.0512248e-07, -1.52033645e-05, -8.576382e-06, 1.5182856e-07, 1.03767775e-07, -1.0871958e-05, -8.732611e-06, 2.6215336e-08, 1.01284385e-07, -6.487446e-06, -8.788768e-06, -9.874178e-08, 9.769532e-08, -2.099805e-06, -8.745291e-06, -2.2164225e-07, 9.303547e-08, 2.2414924e-06, -8.603738e-06, -3.4111443e-07, 8.735144e-08, 6.4880264e-06, -8.366761e-06, -4.5583084e-07, 8.070126e-08, 1.0592969e-05, -8.038073e-06, -5.645231e-07, 7.315401e-08, 1.4511605e-05, -7.6223923e-06, -6.659961e-07, 6.47892e-08, 1.8201816e-05, -7.1253894e-06, -7.591417e-07, 5.5696074e-08, 2.162454e-05, -6.55361e-06, -8.4295095e-07, 4.5972804e-08, 2.4744197e-05, -5.914399e-06, -9.1652595e-07, 3.5725492e-08, 2.7529055e-05, -5.215808e-06, -9.790897e-07, 2.506707e-08, 2.9951567e-05, -4.4665e-06, -1.0299952e-06, 1.4116131e-08, 3.1988646e-05, -3.6756442e-06, -1.0687326e-06, 2.9956015e-09, 3.3621895e-05, -2.8528073e-06, -1.0949349e-06, -8.168631e-09, 3.483778e-05, -2.0078396e-06, -1.1083825e-06, -1.9249171e-08, 3.562773e-05, -1.1507593e-06, -1.1090052e-06, -3.011862e-08, 3.5988207e-05, -2.9163368e-07, -1.0968824e-06, -4.06511e-08, 3.5920697e-05, 5.59538e-07, -1.0722429e-06, -5.0723806e-08, 3.543164e-05, 1.3929415e-06, -1.0354607e-06, -6.021853e-08, 3.453231e-05, 2.199061e-06, -9.870516e-07, -6.902319e-08, 3.3238648e-05, 2.9687892e-06, -9.276652e-07, -7.70332e-08, 3.157102e-05, 3.6935317e-06, -8.5807824e-07, -8.4152944e-08, 2.9553943e-05, 4.365304e-06, -7.7918384e-07, -9.0297e-08, 2.7215754e-05, 4.9768223e-06, -6.919812e-07, -9.53913e-08, 2.458824e-05, 5.521584e-06, -5.9756286e-07, -9.9374176e-08, 2.1706228e-05, 5.9939393e-06, -4.971011e-07, -1.0219725e-07, 1.8607147e-05, 6.3891516e-06, -3.9183377e-07, -1.0382613e-07, 1.533055e-05, 6.703446e-06, -2.8304876e-07, -1.04240975e-07, 1.1917634e-05, 6.9340485e-06, -1.7206814e-07, -1.0343684e-07, 8.410726e-06, 7.079208e-06, -6.023198e-08, -1.0142383e-07, 4.852769e-06, 7.138211e-06, 5.1118253e-08, -9.82271e-08, 1.2868036e-06, 7.111381e-06, 1.6065611e-07, -9.3886534e-08, -2.2445479e-06, 7.0000647e-06, 2.6708645e-07, -8.8456424e-08, -5.6995873e-06, 6.806607e-06, 3.691611e-07, -8.2004725e-08, -9.038031e-06, 6.5343133e-06, 4.656943e-07, -7.4612295e-08, -1.2221478e-05, 6.1874016e-06, 5.555767e-07, -6.6371875e-08, -1.5213853e-05, 5.770941e-06, 6.3778896e-07, -5.738693e-08, -1.7981813e-05, 5.2907844e-06, 7.114137e-07, -4.777032e-08, -2.0495121e-05, 4.7534872e-06, 7.7564624e-07, -3.764284e-08, -2.2726977e-05, 4.1662224e-06, 8.298041e-07, -2.7131675e-08, -2.46543e-05, 3.5366854e-06, 8.7333456e-07, -1.636872e-08, -2.6257969e-05, 2.8729953e-06, 9.058206e-07, -5.48886e-09, -2.7523005e-05, 2.1835913e-06, 9.2698525e-07, 5.3718012e-09, -2.843871e-05, 1.4771254e-06, 9.36694e-07, 1.6077742e-08, -2.8998735e-05, 7.62354e-07, 9.3495527e-07, 2.6495812e-08, -2.9201123e-05, 4.802945e-08, 9.2191925e-07, 3.649699e-08, -2.9048262e-05, -6.572079e-07, 8.978748e-07, 4.595808e-08, -2.8546814e-05, -1.3449348e-06, 8.6324457e-07, 5.4763348e-08, -2.7707574e-05, -2.0070468e-06, 8.185786e-07, 6.2806045e-08, -2.6545295e-05, -2.6358537e-06, 7.64546e-07, 6.998978e-08, -2.5078443e-05, -3.224171e-06, 7.0192544e-07, 7.622982e-08, -2.3328943e-05, -3.765402e-06, 6.315944e-07, 8.1454104e-08, -2.132185e-05, -4.2536126e-06, 5.545168e-07, 8.560424e-08, -1.9085008e-05, -4.683596e-06, 4.717299e-07, 8.8636185e-08, -1.6648668e-05, -5.0509307e-06, 3.843304e-07, 9.052074e-08, -1.404509e-05, -5.3520216e-06, 2.9345995e-07, 9.124394e-08, -1.1308117e-05, -5.5841374e-06, 2.0028985e-07, 9.080708e-08, -8.4727335e-06, -5.7454317e-06, 1.060059e-07, 8.922665e-08, -5.5746254e-06, -5.8349547e-06, 1.1793107e-08, 8.653403e-08, -2.6497305e-06, -5.852653e-06, -8.11795e-08, 8.2774925e-08, 2.662109e-07, -5.7993584e-06, -1.7177365e-07, 7.800867e-08, 3.1380905e-06, -5.6767653e-06, -2.58896e-07, 7.230735e-08, 5.9318554e-06, -5.487397e-06, -3.415116e-07, 6.575468e-08, 8.614915e-06, -5.234563e-06, -4.186564e-07, 5.8444844e-08, 1.1156516e-05, -4.9223067e-06, -4.8944884e-07, 5.048106e-08, 1.35281e-05, -4.555343e-06, -5.530998e-07, 4.197415e-08, 1.570362e-05, -4.1389917e-06, -6.089219e-07, 3.304097e-08, 1.7659822e-05, -3.6790993e-06, -6.5633645e-07, 2.380274e-08, 1.9376495e-05, -3.1819607e-06, -6.948797e-07, 1.4383385e-08, 2.0836665e-05, -2.6542316e-06, -7.2420727e-07, 4.907812e-09, 2.202676e-05, -2.1028407e-06, -7.4409644e-07, -4.4997925e-09, 2.293672e-05, -1.5348982e-06, -7.544476e-07, -1.371764e-08, 2.356007e-05, -9.576042e-07, -7.5528357e-07, -2.2627969e-08, 2.3893934e-05, -3.7815727e-07, -7.467473e-07, -3.1118592e-08, 2.393902e-05, 1.9633609e-07, -7.2909836e-07, -3.908437e-08, 2.3699544e-05, 7.589485e-07, -7.0270767e-07, -4.6428532e-08, 2.3183127e-05, 1.3030154e-06, -6.6805103e-07, -5.3063903e-08, 2.2400638e-05, 1.8222148e-06, -6.257011e-07, -5.8913965e-08, 2.1366006e-05, 2.3106395e-06, -5.763184e-07, -6.3913745e-08, 2.0095997e-05, 2.7628648e-06, -5.2064166e-07, -6.801054e-08, 1.8609955e-05, 3.1740074e-06, -4.5947658e-07, -7.1164486e-08, 1.692952e-05, 3.5397777e-06, -3.936844e-07, -7.334889e-08, 1.5078321e-05, 3.8565217e-06, -3.2416983e-07, -7.455041e-08, 1.3081642e-05, 4.1212575e-06, -2.5186873e-07, -7.476901e-08, 1.09660905e-05, 4.3316973e-06, -1.7773522e-07, -7.401783e-08, 8.759238e-06, 4.486266e-06, -1.027292e-07, -7.23227e-08, 6.4892656e-06, 4.5841057e-06, -2.7803862e-08, -6.9721644e-08, 4.1846015e-06, 4.6250743e-06, 4.610653e-08, -6.626416e-08, 1.873571e-06, 4.6097334e-06, 1.1809828e-07, -6.201031e-08, -4.1595456e-07, 4.5393263e-06, 1.8730934e-07, -5.7029773e-08, -2.6568903e-06, 4.4157523e-06, 2.5292962e-07, -5.140069e-08, -4.8232564e-06, 4.2415263e-06, 3.1421035e-07, -4.5208456e-08, -6.8904765e-06, 4.0197383e-06, 3.7047252e-07, -3.854442e-08, -8.835653e-06, 3.7540026e-06, 4.2111424e-07, -3.150455e-08, -1.0637814e-05, 3.4484015e-06, 4.6561675e-07, -2.4187996e-08, -1.2278134e-05, 3.1074248e-06, 5.035496e-07, -1.669571e-08, -1.3740121e-05, 2.7359067e-06, 5.345741e-07, -9.129019e-09, -1.5009772e-05, 2.3389575e-06, 5.5844583e-07, -1.5882398e-09, -1.6075694e-05, 1.9218949e-06, 5.7501575e-07, 5.8286753e-09, -1.6929189e-05, 1.4901724e-06, 5.8422995e-07, 1.3027422e-08, -1.7564307e-05, 1.0493103e-06, 5.8612835e-07, 1.9918554e-08, -1.797786e-05, 6.048245e-07, 5.8084197e-07, 2.6418604e-08, -1.81694e-05, 1.621589e-07, 5.6858937e-07, 3.2451087e-08, -1.814117e-05, -2.733809e-07, 5.4967154e-07, 3.79474e-08, -1.7898023e-05, -6.9668994e-07, 5.2446654e-07, 4.2847574e-08, -1.7447295e-05, -1.1029227e-06, 4.934227e-07, 4.7100894e-08, -1.6798671e-05, -1.4875471e-06, 4.5705104e-07, 5.066639e-08, -1.5964017e-05, -1.8463934e-06, 4.159176e-07, 5.3513162e-08, -1.4957177e-05, -2.175697e-06, 3.7063478e-07, 5.562056e-08, -1.3793775e-05, -2.4721362e-06, 3.2185224e-07, 5.6978227e-08, -1.2490975e-05, -2.7328622e-06, 2.7024802e-07, 5.7585982e-08, -1.1067243e-05, -2.955523e-06, 2.1651901e-07, 5.745359e-08, -9.542092e-06, -3.1382815e-06, 1.6137176e-07, 5.6600356e-08, -7.935824e-06, -3.2798243e-06, 1.0551322e-07, 5.505465e-08, -6.2692657e-06, -3.3793672e-06, 4.964183e-08, 5.2853252e-08, -4.5635034e-06, -3.4366499e-06, -5.5610947e-09, 5.0040686e-08, -2.8396234e-06, -3.4519285e-06, -5.943951e-08, 4.6668365e-08, -1.1184601e-06, -3.4259588e-06, -1.1137024e-07, 4.2793744e-08, 5.796517e-07, -3.3599742e-06, -1.6076991e-07, 3.847936e-08, 2.235108e-06, -3.255661e-06, -2.0710128e-07, 3.379185e-08, 3.8292546e-06, -3.1151246e-06, -2.498786e-07, 2.8800953e-08, 5.3445865e-06, -2.940854e-06, -2.886724e-07, 2.357846e-08, 6.764932e-06, -2.7356832e-06, -3.2311326e-07, 1.8197206e-08, 8.075614e-06, -2.5027464e-06, -3.528947e-07, 1.2730045e-08, 9.263586e-06, -2.2454342e-06, -3.7777525e-07, 7.2488784e-09, 1.0317554e-05, -1.9673455e-06, -3.9757973e-07, 1.8237177e-09, 1.1228064e-05, -1.6722387e-06, -4.1219926e-07, -3.478203e-09, 1.198757e-05, -1.3639828e-06, -4.2159098e-07, -8.59324e-09, 1.2590479e-05, -1.0465085e-06, -4.2577645e-07, -1.34620795e-08, 1.3033169e-05, -7.237587e-07, -4.248397e-07, -1.8030399e-08, 1.3313982e-05, -3.996422e-07, -4.189241e-07, -2.2249425e-08, 1.3433195e-05, -7.798749e-08, -4.0822906e-07, -2.6076421e-08, 1.33929725e-05, 2.3750053e-07, -3.9300585e-07, -2.9475036e-08, 1.319729e-05, 5.4328103e-07, -3.7355287e-07, -3.2415596e-08, 1.2851847e-05, 8.360148e-07, -3.5021077e-07, -3.4875267e-08, 1.2363951e-05, 1.1125984e-06, -3.2335683e-07, -3.683812e-08, 1.17424e-05, 1.3701942e-06, -2.9339944e-07, -3.8295113e-08, 1.0997336e-05, 1.6062565e-06, -2.6077205e-07, -3.9243965e-08, 1.0140098e-05, 1.8185539e-06, -2.2592734e-07, -3.968895e-08, 9.183057e-06, 2.005186e-06, -1.89331e-07, -3.9640597e-08, 8.13945e-06, 2.1645976e-06, -1.5145595e-07, -3.911534e-08, 7.0232013e-06, 2.2955874e-06, -1.1277631e-07, -3.8135074e-08, 5.848748e-06, 2.3973107e-06, -7.376182e-08, -3.6726675e-08, 4.63086e-06, 2.4692815e-06, -3.487238e-08, -3.492145e-08, 3.384461e-06, 2.5113677e-06, 3.4470127e-09, -3.275457e-08, 2.124454e-06, 2.523782e-06, 4.077105e-08, -3.0264463e-08, 8.655517e-07, 2.5070717e-06, 7.6698434e-08, -2.7492183e-08, -3.7788712e-07, 2.4621015e-06, 1.1085578e-07, -2.4480785e-08, -1.5920119e-06, 2.3900368e-06, 1.4290102e-07, -2.1274682e-08, -2.7636254e-06, 2.292321e-06, 1.7252636e-07, -1.7919024e-08, -3.8803164e-06, 2.170652e-06, 1.9946066e-07, -1.4459092e-08, -4.930582e-06, 2.0269558e-06, 2.2347136e-07, -1.09397105e-08, -5.903931e-06, 1.8633597e-06, 2.4436585e-07, -7.404702e-09, -6.790983e-06, 1.6821613e-06, 2.619923e-07, -3.896372e-09, -7.5835414e-06, 1.4857994e-06, 2.7624012e-07, -4.5504253e-10, -8.274657e-06, 1.2768228e-06, 2.8703965e-07, 2.8813676e-09, -8.8586785e-06, 1.0578584e-06, 2.9436183e-07, 6.0777094e-09, -9.331277e-06, 8.315807e-07, 2.9821695e-07, 9.101918e-09, -9.689472e-06, 6.0068055e-07, 2.9865333e-07, 1.1925269e-08, -9.9316185e-06, 3.6783518e-07, 2.9575557e-07, 1.4522579e-08, -1.0057409e-05, 1.3567924e-07, 2.8964226e-07, 1.687235e-08, -1.006783e-05, -9.3223015e-08, 2.804638e-07, 1.895686e-08, -9.9651315e-06, -3.1640386e-07, 2.683995e-07, 2.076219e-08, -9.752765e-06, -5.315164e-07, 2.5365483e-07, 2.2278224e-08, -9.4353245e-06, -7.363568e-07, 2.364583e-07, 2.3498568e-08, -9.018461e-06, -9.2888484e-07, 2.1705834e-07, 2.4420462e-08, -8.508804e-06, -1.1072412e-06, 1.9571996e-07, 2.504461e-08, -7.913864e-06, -1.2697633e-06, 1.7272144e-07, 2.5375021e-08, -7.241929e-06, -1.414998e-06, 1.4835106e-07, 2.541878e-08, -6.5019617e-06, -1.541712e-06, 1.2290369e-07, 2.5185816e-08, -5.7034827e-06, -1.6488997e-06, 9.667761e-08, 2.4688644e-08, -4.856458e-06, -1.7357884e-06, 6.9971286e-08, 2.394209e-08, -3.971181e-06, -1.8018407e-06, 4.308036e-08, 2.2962999e-08, -3.0581555e-06, -1.8467547e-06, 1.629469e-08, 2.1769953e-08, -2.127977e-06, -1.870462e-06, -1.0104367e-08, 2.0382977e-08, -1.191218e-06, -1.8731229e-06, -3.584656e-08, 1.8823236e-08, -2.5831505e-07, -1.8551193e-06, -6.0675106e-08, 1.7112768e-08, 6.6053957e-07, -1.8170463e-06, -8.4348855e-08, 1.527419e-08, 1.5555025e-06, -1.7597008e-06, -1.0664425e-07, 1.3330456e-08, 2.4171766e-06, -1.6840693e-06, -1.2735704e-07, 1.1304585e-08, 3.2367025e-06, -1.5913134e-06, -1.4630375e-07, 9.219448e-09, 4.005842e-06, -1.4827542e-06, -1.6332292e-07, 7.0975457e-09, 4.717054e-06, -1.3598553e-06, -1.7827617e-07, 4.9608166e-09, 5.3635604e-06, -1.2242051e-06, -1.9104887e-07, 2.830462e-09, 5.9394056e-06, -1.0774975e-06, -2.0155073e-07, 7.267915e-10, 6.4395026e-06, -9.2151265e-07, -2.097161e-07, -1.3309103e-09, 6.859673e-06, -7.5809737e-07, -2.1550403e-07, -3.3244987e-09, 7.196672e-06, -5.8914435e-07, -2.1889811e-07, -5.237066e-09, 7.4482105e-06, -4.1657208e-07, -2.1990613e-07, -7.0530164e-09, 7.6129595e-06, -2.423047e-07, -2.1855952e-07, -8.758133e-09, 7.690551e-06, -6.825226e-08, -2.1491257e-07, -1.0339618e-08, 7.681562e-06, 1.0370888e-07, -2.0904156e-07, -1.1786129e-08, 7.5874973e-06, 2.7175466e-07, -2.0104353e-07, -1.30878e-08, 7.4107566e-06, 4.3413118e-07, -1.9103518e-07, -1.4236247e-08, 7.1545946e-06, 5.891718e-07, -1.7915134e-07, -1.522457e-08, 6.8230747e-06, 7.353128e-07, -1.6554344e-07, -1.6047345e-08, 6.421014e-06, 8.7110806e-07, -1.5037789e-07, -1.670061e-08, 5.953919e-06, 9.952423e-07, -1.3383429e-07, -1.7181845e-08, 5.42792e-06, 1.1065426e-06, -1.1610354e-07, -1.7489937e-08, 4.8496945e-06, 1.2039893e-06, -9.738596e-08, -1.7625162e-08, 4.2263923e-06, 1.2867233e-06, -7.7889204e-08, -1.7589148e-08, 3.5655482e-06, 1.3540545e-06, -5.7826295e-08, -1.7384838e-08, 2.875001e-06, 1.4054654e-06, -3.741348e-08, -1.7016449e-08, 2.1628027e-06, 1.4406153e-06, -1.6868164e-08, -1.648943e-08, 1.4371319e-06, 1.4593417e-06, 3.5931949e-09, -1.5810418e-08, 7.0620405e-07, 1.46166e-06, 2.3757162e-08, -1.4987192e-08, -2.181738e-08, 1.447761e-06, 4.3415373e-08, -1.4028609e-08, -7.389075e-07, 1.4180075e-06, 6.236653e-08, -1.2944563e-08, -1.4372646e-06, 1.3729289e-06, 8.0418324e-08, -1.1745907e-08, -2.1093917e-06, 1.3132131e-06, 9.7389275e-08, -1.0444398e-08, -2.7481738e-06, 1.2396989e-06, 1.1311048e-07, -9.0526155e-09};
endpackage
`endif
