`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam N = 4;
	localparam M = 4;
	localparam real Lfr[0:3] = {0.923863, 0.923863, 0.8888867, 0.8888867};
	localparam real Lfi[0:3] = {0.22634004, -0.22634004, 0.0844262, -0.0844262};
	localparam real Lbr[0:3] = {0.923863, 0.923863, 0.8888867, 0.8888867};
	localparam real Lbi[0:3] = {0.22634004, -0.22634004, 0.0844262, -0.0844262};
	localparam real Wfr[0:3] = {0.007497563, 0.007497563, -0.0020543877, -0.0020543877};
	localparam real Wfi[0:3] = {0.0014516033, -0.0014516033, -0.0048014303, 0.0048014303};
	localparam real Wbr[0:3] = {-0.007497563, -0.007497563, 0.0020543877, 0.0020543877};
	localparam real Wbi[0:3] = {-0.0014516033, 0.0014516033, 0.0048014303, -0.0048014303};
	localparam real Ffr[0:3][0:99] = '{
		'{1.5881557, 0.7547344, -0.42185825, 0.007546211, 1.8962913, 0.48151, -0.42255256, 0.038024865, 2.0669386, 0.2068506, -0.39908394, 0.063432075, 2.1034615, -0.053444244, -0.35509223, 0.082802005, 2.0165524, -0.28589895, -0.2950409, 0.095605075, 1.822924, -0.47990912, -0.2238841, 0.10173665, 1.5437828, -0.62807274, -0.14673743, 0.10148251, 1.2031924, -0.7263073, -0.06857083, 0.09546536, 0.82642823, -0.7737664, 0.006060983, 0.08457727, 0.43842137, -0.7725798, 0.07323868, 0.069903076, 0.062369436, -0.72744864, 0.12984131, 0.05264022, -0.2814213, -0.64513206, 0.1736483, 0.03401971, -0.57641834, -0.5338663, 0.2033802, 0.015232723, -0.81044656, -0.4027536, 0.21868213, -0.0026335253, -0.9759671, -0.2611614, 0.22005586, -0.018647881, -1.0700662, -0.11816227, 0.20874971, -0.032073487, -1.0941802, 0.017954962, 0.18661615, -0.042391293, -1.0536001, 0.14008348, 0.15594865, -0.049308926, -0.9568018, 0.2425911, 0.11930892, -0.052755747, -0.8146601, 0.321501, 0.07935524, -0.052865785, -0.6395996, 0.37456077, 0.038681667, -0.049950585, -0.44473895, 0.40120682, -0.0003237382, -0.044464532, -0.2430763, 0.40243542, -0.035595525, -0.03696535, -0.046759624, 0.38059747, -0.06547787, -0.028072434, 0.13352495, 0.33913532, -0.08878002, -0.018425668},
		'{1.5881557, 0.7547344, -0.42185825, 0.007546211, 1.8962913, 0.48151, -0.42255256, 0.038024865, 2.0669386, 0.2068506, -0.39908394, 0.063432075, 2.1034615, -0.053444244, -0.35509223, 0.082802005, 2.0165524, -0.28589895, -0.2950409, 0.095605075, 1.822924, -0.47990912, -0.2238841, 0.10173665, 1.5437828, -0.62807274, -0.14673743, 0.10148251, 1.2031924, -0.7263073, -0.06857083, 0.09546536, 0.82642823, -0.7737664, 0.006060983, 0.08457727, 0.43842137, -0.7725798, 0.07323868, 0.069903076, 0.062369436, -0.72744864, 0.12984131, 0.05264022, -0.2814213, -0.64513206, 0.1736483, 0.03401971, -0.57641834, -0.5338663, 0.2033802, 0.015232723, -0.81044656, -0.4027536, 0.21868213, -0.0026335253, -0.9759671, -0.2611614, 0.22005586, -0.018647881, -1.0700662, -0.11816227, 0.20874971, -0.032073487, -1.0941802, 0.017954962, 0.18661615, -0.042391293, -1.0536001, 0.14008348, 0.15594865, -0.049308926, -0.9568018, 0.2425911, 0.11930892, -0.052755747, -0.8146601, 0.321501, 0.07935524, -0.052865785, -0.6395996, 0.37456077, 0.038681667, -0.049950585, -0.44473895, 0.40120682, -0.0003237382, -0.044464532, -0.2430763, 0.40243542, -0.035595525, -0.03696535, -0.046759624, 0.38059747, -0.06547787, -0.028072434, 0.13352495, 0.33913532, -0.08878002, -0.018425668},
		'{-1.3553582, -0.65067863, 0.3077727, -0.2458136, -1.6303499, -0.46066287, 0.22754894, -0.20613672, -1.8178369, -0.3002024, 0.15915948, -0.17049015, -1.9319099, -0.1664296, 0.10153671, -0.1387509, -1.9852324, -0.056538545, 0.053619795, -0.110744834, -1.9890833, 0.032172833, 0.014373968, -0.08626044, -1.953418, 0.10227121, -0.01719458, -0.06506049, -1.8869433, 0.15616533, -0.042027675, -0.046891894, -1.7972002, 0.19609112, -0.061007347, -0.031493865, -1.6906543, 0.22410317, -0.074950784, -0.018604517, -1.572787, 0.24207154, -0.084607564, -0.007966216, -1.4481893, 0.25168267, -0.09065877, 0.00067027594, -1.3206521, 0.25444388, -0.09371758, 0.0075426428, -1.1932551, 0.2516902, -0.09433117, 0.012874734, -1.0684508, 0.24459344, -0.09298334, 0.016875006, -0.94814396, 0.23417237, -0.09009804, 0.019735591, -0.83376557, 0.22130394, -0.08604318, 0.021631854, -0.72634095, 0.20673496, -0.08113485, 0.022722388, -0.6265522, 0.19109392, -0.07564168, 0.023149317, -0.5347945, 0.1749028, -0.06978922, 0.023038877, -0.45122632, 0.15858841, -0.0637643, 0.02250217, -0.37581468, 0.14249347, -0.057719193, 0.021636076, -0.30837435, 0.12688692, -0.05177573, 0.020524247, -0.24860243, 0.111973636, -0.046029046, 0.019238153, -0.19610818, 0.0979035, -0.04055115, 0.017838178},
		'{-1.3553582, -0.65067863, 0.3077727, -0.2458136, -1.6303499, -0.46066287, 0.22754894, -0.20613672, -1.8178369, -0.3002024, 0.15915948, -0.17049015, -1.9319099, -0.1664296, 0.10153671, -0.1387509, -1.9852324, -0.056538545, 0.053619795, -0.110744834, -1.9890833, 0.032172833, 0.014373968, -0.08626044, -1.953418, 0.10227121, -0.01719458, -0.06506049, -1.8869433, 0.15616533, -0.042027675, -0.046891894, -1.7972002, 0.19609112, -0.061007347, -0.031493865, -1.6906543, 0.22410317, -0.074950784, -0.018604517, -1.572787, 0.24207154, -0.084607564, -0.007966216, -1.4481893, 0.25168267, -0.09065877, 0.00067027594, -1.3206521, 0.25444388, -0.09371758, 0.0075426428, -1.1932551, 0.2516902, -0.09433117, 0.012874734, -1.0684508, 0.24459344, -0.09298334, 0.016875006, -0.94814396, 0.23417237, -0.09009804, 0.019735591, -0.83376557, 0.22130394, -0.08604318, 0.021631854, -0.72634095, 0.20673496, -0.08113485, 0.022722388, -0.6265522, 0.19109392, -0.07564168, 0.023149317, -0.5347945, 0.1749028, -0.06978922, 0.023038877, -0.45122632, 0.15858841, -0.0637643, 0.02250217, -0.37581468, 0.14249347, -0.057719193, 0.021636076, -0.30837435, 0.12688692, -0.05177573, 0.020524247, -0.24860243, 0.111973636, -0.046029046, 0.019238153, -0.19610818, 0.0979035, -0.04055115, 0.017838178}};
	localparam real Ffi[0:3][0:99] = '{
		'{-1.895612, 0.9532613, 0.14497346, -0.1371971, -1.3918226, 1.0515095, 0.038452197, -0.12504332, -0.8566468, 1.0804358, -0.060116, -0.10691635, -0.32359335, 1.0449932, -0.14586763, -0.08441885, 0.17714167, 0.953334, -0.2151333, -0.05925004, 0.6200812, 0.8160396, -0.26553327, -0.033099666, 0.9854708, 0.6452862, -0.29599032, -0.00755248, 1.2598599, 0.45399803, -0.30666706, 0.0159921, 1.4362686, 0.25503957, -0.29883868, 0.036382142, 1.5139693, 0.06048731, -0.27471414, 0.05275534, 1.4979326, -0.11898376, -0.2372214, 0.06456057, 1.3980012, -0.27457544, -0.1897718, 0.07155971, 1.2278646, -0.39968932, -0.13601959, 0.0738114, 1.0039122, -0.4900935, -0.079630375, 0.071639396, 0.74404085, -0.5439385, -0.024071041, 0.065588914, 0.46649137, -0.561636, 0.02756911, 0.056374412, 0.18877532, -0.54561955, 0.0727185, 0.04482272, -0.07325427, -0.5000138, 0.10942064, 0.03181521, -0.3061488, -0.43023777, 0.13638711, 0.018232308, -0.4994021, -0.3425727, 0.15300739, 0.0049034175, -0.64576936, -0.2437217, 0.15931915, -0.007435558, -0.7413694, -0.14038736, 0.15594427, -0.018175256, -0.785586, -0.038889512, 0.14399788, -0.02685555, -0.78079176, 0.05515867, 0.12497762, -0.033177588, -0.7319282, 0.1371035, 0.100641936, -0.03700546},
		'{1.895612, -0.9532613, -0.14497346, 0.1371971, 1.3918226, -1.0515095, -0.038452197, 0.12504332, 0.8566468, -1.0804358, 0.060116, 0.10691635, 0.32359335, -1.0449932, 0.14586763, 0.08441885, -0.17714167, -0.953334, 0.2151333, 0.05925004, -0.6200812, -0.8160396, 0.26553327, 0.033099666, -0.9854708, -0.6452862, 0.29599032, 0.00755248, -1.2598599, -0.45399803, 0.30666706, -0.0159921, -1.4362686, -0.25503957, 0.29883868, -0.036382142, -1.5139693, -0.06048731, 0.27471414, -0.05275534, -1.4979326, 0.11898376, 0.2372214, -0.06456057, -1.3980012, 0.27457544, 0.1897718, -0.07155971, -1.2278646, 0.39968932, 0.13601959, -0.0738114, -1.0039122, 0.4900935, 0.079630375, -0.071639396, -0.74404085, 0.5439385, 0.024071041, -0.065588914, -0.46649137, 0.561636, -0.02756911, -0.056374412, -0.18877532, 0.54561955, -0.0727185, -0.04482272, 0.07325427, 0.5000138, -0.10942064, -0.03181521, 0.3061488, 0.43023777, -0.13638711, -0.018232308, 0.4994021, 0.3425727, -0.15300739, -0.0049034175, 0.64576936, 0.2437217, -0.15931915, 0.007435558, 0.7413694, 0.14038736, -0.15594427, 0.018175256, 0.785586, 0.038889512, -0.14399788, 0.02685555, 0.78079176, -0.05515867, -0.12497762, 0.033177588, 0.7319282, -0.1371035, -0.100641936, 0.03700546},
		'{5.0409703, -1.3943145, 0.5451638, -0.14644392, 4.3664236, -1.294322, 0.5105729, -0.15092516, 3.7436113, -1.1893976, 0.47305256, -0.15155871, 3.1741734, -1.0825846, 0.43392736, -0.14911234, 2.6583765, -0.9763461, 0.3942846, -0.1442582, 2.19539, -0.87263435, 0.35500127, -0.13757895, 1.7835221, -0.77295685, 0.31676942, -0.12957475, 1.4204293, -0.6784367, 0.28012046, -0.12067007, 1.1032933, -0.5898689, 0.24544711, -0.111220926, 0.8289719, -0.5077714, 0.21302405, -0.10152171, 0.5941266, -0.43243104, 0.18302643, -0.091812, 0.3953268, -0.363945, 0.15554667, -0.08228303, 0.2291356, -0.30225727, 0.13060938, -0.0730837, 0.09217794, -0.24719071, 0.10818472, -0.06432633, -0.018806256, -0.19847529, 0.088199936, -0.056091852, -0.106921874, -0.15577194, 0.07054952, -0.048434608, -0.17508963, -0.11869333, 0.05510389, -0.041386675, -0.22602649, -0.086821064, 0.041716818, -0.03496177, -0.26223415, -0.059720244, 0.030231616, -0.029158687, -0.28599387, -0.036951195, 0.02048634, -0.02396436, -0.2993668, -0.018079046, 0.0123179965, -0.019356515, -0.3041985, -0.0026812062, 0.005565926, -0.015305976, -0.30212662, 0.009646894, 7.446508e-05, -0.011778627, -0.2945912, 0.019287577, -0.0043050377, -0.00873708, -0.28284675, 0.026597979, -0.007712748, -0.00614207},
		'{-5.0409703, 1.3943145, -0.5451638, 0.14644392, -4.3664236, 1.294322, -0.5105729, 0.15092516, -3.7436113, 1.1893976, -0.47305256, 0.15155871, -3.1741734, 1.0825846, -0.43392736, 0.14911234, -2.6583765, 0.9763461, -0.3942846, 0.1442582, -2.19539, 0.87263435, -0.35500127, 0.13757895, -1.7835221, 0.77295685, -0.31676942, 0.12957475, -1.4204293, 0.6784367, -0.28012046, 0.12067007, -1.1032933, 0.5898689, -0.24544711, 0.111220926, -0.8289719, 0.5077714, -0.21302405, 0.10152171, -0.5941266, 0.43243104, -0.18302643, 0.091812, -0.3953268, 0.363945, -0.15554667, 0.08228303, -0.2291356, 0.30225727, -0.13060938, 0.0730837, -0.09217794, 0.24719071, -0.10818472, 0.06432633, 0.018806256, 0.19847529, -0.088199936, 0.056091852, 0.106921874, 0.15577194, -0.07054952, 0.048434608, 0.17508963, 0.11869333, -0.05510389, 0.041386675, 0.22602649, 0.086821064, -0.041716818, 0.03496177, 0.26223415, 0.059720244, -0.030231616, 0.029158687, 0.28599387, 0.036951195, -0.02048634, 0.02396436, 0.2993668, 0.018079046, -0.0123179965, 0.019356515, 0.3041985, 0.0026812062, -0.005565926, 0.015305976, 0.30212662, -0.009646894, -7.446508e-05, 0.011778627, 0.2945912, -0.019287577, 0.0043050377, 0.00873708, 0.28284675, -0.026597979, 0.007712748, 0.00614207}};
	localparam real Fbr[0:3][0:99] = '{
		'{-1.5881557, 0.7547344, 0.42185825, 0.007546211, -1.8962913, 0.48151, 0.42255256, 0.038024865, -2.0669386, 0.2068506, 0.39908394, 0.063432075, -2.1034615, -0.053444244, 0.35509223, 0.082802005, -2.0165524, -0.28589895, 0.2950409, 0.095605075, -1.822924, -0.47990912, 0.2238841, 0.10173665, -1.5437828, -0.62807274, 0.14673743, 0.10148251, -1.2031924, -0.7263073, 0.06857083, 0.09546536, -0.82642823, -0.7737664, -0.006060983, 0.08457727, -0.43842137, -0.7725798, -0.07323868, 0.069903076, -0.062369436, -0.72744864, -0.12984131, 0.05264022, 0.2814213, -0.64513206, -0.1736483, 0.03401971, 0.57641834, -0.5338663, -0.2033802, 0.015232723, 0.81044656, -0.4027536, -0.21868213, -0.0026335253, 0.9759671, -0.2611614, -0.22005586, -0.018647881, 1.0700662, -0.11816227, -0.20874971, -0.032073487, 1.0941802, 0.017954962, -0.18661615, -0.042391293, 1.0536001, 0.14008348, -0.15594865, -0.049308926, 0.9568018, 0.2425911, -0.11930892, -0.052755747, 0.8146601, 0.321501, -0.07935524, -0.052865785, 0.6395996, 0.37456077, -0.038681667, -0.049950585, 0.44473895, 0.40120682, 0.0003237382, -0.044464532, 0.2430763, 0.40243542, 0.035595525, -0.03696535, 0.046759624, 0.38059747, 0.06547787, -0.028072434, -0.13352495, 0.33913532, 0.08878002, -0.018425668},
		'{-1.5881557, 0.7547344, 0.42185825, 0.007546211, -1.8962913, 0.48151, 0.42255256, 0.038024865, -2.0669386, 0.2068506, 0.39908394, 0.063432075, -2.1034615, -0.053444244, 0.35509223, 0.082802005, -2.0165524, -0.28589895, 0.2950409, 0.095605075, -1.822924, -0.47990912, 0.2238841, 0.10173665, -1.5437828, -0.62807274, 0.14673743, 0.10148251, -1.2031924, -0.7263073, 0.06857083, 0.09546536, -0.82642823, -0.7737664, -0.006060983, 0.08457727, -0.43842137, -0.7725798, -0.07323868, 0.069903076, -0.062369436, -0.72744864, -0.12984131, 0.05264022, 0.2814213, -0.64513206, -0.1736483, 0.03401971, 0.57641834, -0.5338663, -0.2033802, 0.015232723, 0.81044656, -0.4027536, -0.21868213, -0.0026335253, 0.9759671, -0.2611614, -0.22005586, -0.018647881, 1.0700662, -0.11816227, -0.20874971, -0.032073487, 1.0941802, 0.017954962, -0.18661615, -0.042391293, 1.0536001, 0.14008348, -0.15594865, -0.049308926, 0.9568018, 0.2425911, -0.11930892, -0.052755747, 0.8146601, 0.321501, -0.07935524, -0.052865785, 0.6395996, 0.37456077, -0.038681667, -0.049950585, 0.44473895, 0.40120682, 0.0003237382, -0.044464532, 0.2430763, 0.40243542, 0.035595525, -0.03696535, 0.046759624, 0.38059747, 0.06547787, -0.028072434, -0.13352495, 0.33913532, 0.08878002, -0.018425668},
		'{1.3553582, -0.65067863, -0.3077727, -0.2458136, 1.6303499, -0.46066287, -0.22754894, -0.20613672, 1.8178369, -0.3002024, -0.15915948, -0.17049015, 1.9319099, -0.1664296, -0.10153671, -0.1387509, 1.9852324, -0.056538545, -0.053619795, -0.110744834, 1.9890833, 0.032172833, -0.014373968, -0.08626044, 1.953418, 0.10227121, 0.01719458, -0.06506049, 1.8869433, 0.15616533, 0.042027675, -0.046891894, 1.7972002, 0.19609112, 0.061007347, -0.031493865, 1.6906543, 0.22410317, 0.074950784, -0.018604517, 1.572787, 0.24207154, 0.084607564, -0.007966216, 1.4481893, 0.25168267, 0.09065877, 0.00067027594, 1.3206521, 0.25444388, 0.09371758, 0.0075426428, 1.1932551, 0.2516902, 0.09433117, 0.012874734, 1.0684508, 0.24459344, 0.09298334, 0.016875006, 0.94814396, 0.23417237, 0.09009804, 0.019735591, 0.83376557, 0.22130394, 0.08604318, 0.021631854, 0.72634095, 0.20673496, 0.08113485, 0.022722388, 0.6265522, 0.19109392, 0.07564168, 0.023149317, 0.5347945, 0.1749028, 0.06978922, 0.023038877, 0.45122632, 0.15858841, 0.0637643, 0.02250217, 0.37581468, 0.14249347, 0.057719193, 0.021636076, 0.30837435, 0.12688692, 0.05177573, 0.020524247, 0.24860243, 0.111973636, 0.046029046, 0.019238153, 0.19610818, 0.0979035, 0.04055115, 0.017838178},
		'{1.3553582, -0.65067863, -0.3077727, -0.2458136, 1.6303499, -0.46066287, -0.22754894, -0.20613672, 1.8178369, -0.3002024, -0.15915948, -0.17049015, 1.9319099, -0.1664296, -0.10153671, -0.1387509, 1.9852324, -0.056538545, -0.053619795, -0.110744834, 1.9890833, 0.032172833, -0.014373968, -0.08626044, 1.953418, 0.10227121, 0.01719458, -0.06506049, 1.8869433, 0.15616533, 0.042027675, -0.046891894, 1.7972002, 0.19609112, 0.061007347, -0.031493865, 1.6906543, 0.22410317, 0.074950784, -0.018604517, 1.572787, 0.24207154, 0.084607564, -0.007966216, 1.4481893, 0.25168267, 0.09065877, 0.00067027594, 1.3206521, 0.25444388, 0.09371758, 0.0075426428, 1.1932551, 0.2516902, 0.09433117, 0.012874734, 1.0684508, 0.24459344, 0.09298334, 0.016875006, 0.94814396, 0.23417237, 0.09009804, 0.019735591, 0.83376557, 0.22130394, 0.08604318, 0.021631854, 0.72634095, 0.20673496, 0.08113485, 0.022722388, 0.6265522, 0.19109392, 0.07564168, 0.023149317, 0.5347945, 0.1749028, 0.06978922, 0.023038877, 0.45122632, 0.15858841, 0.0637643, 0.02250217, 0.37581468, 0.14249347, 0.057719193, 0.021636076, 0.30837435, 0.12688692, 0.05177573, 0.020524247, 0.24860243, 0.111973636, 0.046029046, 0.019238153, 0.19610818, 0.0979035, 0.04055115, 0.017838178}};
	localparam real Fbi[0:3][0:99] = '{
		'{1.895612, 0.9532613, -0.14497346, -0.1371971, 1.3918226, 1.0515095, -0.038452197, -0.12504332, 0.8566468, 1.0804358, 0.060116, -0.10691635, 0.32359335, 1.0449932, 0.14586763, -0.08441885, -0.17714167, 0.953334, 0.2151333, -0.05925004, -0.6200812, 0.8160396, 0.26553327, -0.033099666, -0.9854708, 0.6452862, 0.29599032, -0.00755248, -1.2598599, 0.45399803, 0.30666706, 0.0159921, -1.4362686, 0.25503957, 0.29883868, 0.036382142, -1.5139693, 0.06048731, 0.27471414, 0.05275534, -1.4979326, -0.11898376, 0.2372214, 0.06456057, -1.3980012, -0.27457544, 0.1897718, 0.07155971, -1.2278646, -0.39968932, 0.13601959, 0.0738114, -1.0039122, -0.4900935, 0.079630375, 0.071639396, -0.74404085, -0.5439385, 0.024071041, 0.065588914, -0.46649137, -0.561636, -0.02756911, 0.056374412, -0.18877532, -0.54561955, -0.0727185, 0.04482272, 0.07325427, -0.5000138, -0.10942064, 0.03181521, 0.3061488, -0.43023777, -0.13638711, 0.018232308, 0.4994021, -0.3425727, -0.15300739, 0.0049034175, 0.64576936, -0.2437217, -0.15931915, -0.007435558, 0.7413694, -0.14038736, -0.15594427, -0.018175256, 0.785586, -0.038889512, -0.14399788, -0.02685555, 0.78079176, 0.05515867, -0.12497762, -0.033177588, 0.7319282, 0.1371035, -0.100641936, -0.03700546},
		'{-1.895612, -0.9532613, 0.14497346, 0.1371971, -1.3918226, -1.0515095, 0.038452197, 0.12504332, -0.8566468, -1.0804358, -0.060116, 0.10691635, -0.32359335, -1.0449932, -0.14586763, 0.08441885, 0.17714167, -0.953334, -0.2151333, 0.05925004, 0.6200812, -0.8160396, -0.26553327, 0.033099666, 0.9854708, -0.6452862, -0.29599032, 0.00755248, 1.2598599, -0.45399803, -0.30666706, -0.0159921, 1.4362686, -0.25503957, -0.29883868, -0.036382142, 1.5139693, -0.06048731, -0.27471414, -0.05275534, 1.4979326, 0.11898376, -0.2372214, -0.06456057, 1.3980012, 0.27457544, -0.1897718, -0.07155971, 1.2278646, 0.39968932, -0.13601959, -0.0738114, 1.0039122, 0.4900935, -0.079630375, -0.071639396, 0.74404085, 0.5439385, -0.024071041, -0.065588914, 0.46649137, 0.561636, 0.02756911, -0.056374412, 0.18877532, 0.54561955, 0.0727185, -0.04482272, -0.07325427, 0.5000138, 0.10942064, -0.03181521, -0.3061488, 0.43023777, 0.13638711, -0.018232308, -0.4994021, 0.3425727, 0.15300739, -0.0049034175, -0.64576936, 0.2437217, 0.15931915, 0.007435558, -0.7413694, 0.14038736, 0.15594427, 0.018175256, -0.785586, 0.038889512, 0.14399788, 0.02685555, -0.78079176, -0.05515867, 0.12497762, 0.033177588, -0.7319282, -0.1371035, 0.100641936, 0.03700546},
		'{-5.0409703, -1.3943145, -0.5451638, -0.14644392, -4.3664236, -1.294322, -0.5105729, -0.15092516, -3.7436113, -1.1893976, -0.47305256, -0.15155871, -3.1741734, -1.0825846, -0.43392736, -0.14911234, -2.6583765, -0.9763461, -0.3942846, -0.1442582, -2.19539, -0.87263435, -0.35500127, -0.13757895, -1.7835221, -0.77295685, -0.31676942, -0.12957475, -1.4204293, -0.6784367, -0.28012046, -0.12067007, -1.1032933, -0.5898689, -0.24544711, -0.111220926, -0.8289719, -0.5077714, -0.21302405, -0.10152171, -0.5941266, -0.43243104, -0.18302643, -0.091812, -0.3953268, -0.363945, -0.15554667, -0.08228303, -0.2291356, -0.30225727, -0.13060938, -0.0730837, -0.09217794, -0.24719071, -0.10818472, -0.06432633, 0.018806256, -0.19847529, -0.088199936, -0.056091852, 0.106921874, -0.15577194, -0.07054952, -0.048434608, 0.17508963, -0.11869333, -0.05510389, -0.041386675, 0.22602649, -0.086821064, -0.041716818, -0.03496177, 0.26223415, -0.059720244, -0.030231616, -0.029158687, 0.28599387, -0.036951195, -0.02048634, -0.02396436, 0.2993668, -0.018079046, -0.0123179965, -0.019356515, 0.3041985, -0.0026812062, -0.005565926, -0.015305976, 0.30212662, 0.009646894, -7.446508e-05, -0.011778627, 0.2945912, 0.019287577, 0.0043050377, -0.00873708, 0.28284675, 0.026597979, 0.007712748, -0.00614207},
		'{5.0409703, 1.3943145, 0.5451638, 0.14644392, 4.3664236, 1.294322, 0.5105729, 0.15092516, 3.7436113, 1.1893976, 0.47305256, 0.15155871, 3.1741734, 1.0825846, 0.43392736, 0.14911234, 2.6583765, 0.9763461, 0.3942846, 0.1442582, 2.19539, 0.87263435, 0.35500127, 0.13757895, 1.7835221, 0.77295685, 0.31676942, 0.12957475, 1.4204293, 0.6784367, 0.28012046, 0.12067007, 1.1032933, 0.5898689, 0.24544711, 0.111220926, 0.8289719, 0.5077714, 0.21302405, 0.10152171, 0.5941266, 0.43243104, 0.18302643, 0.091812, 0.3953268, 0.363945, 0.15554667, 0.08228303, 0.2291356, 0.30225727, 0.13060938, 0.0730837, 0.09217794, 0.24719071, 0.10818472, 0.06432633, -0.018806256, 0.19847529, 0.088199936, 0.056091852, -0.106921874, 0.15577194, 0.07054952, 0.048434608, -0.17508963, 0.11869333, 0.05510389, 0.041386675, -0.22602649, 0.086821064, 0.041716818, 0.03496177, -0.26223415, 0.059720244, 0.030231616, 0.029158687, -0.28599387, 0.036951195, 0.02048634, 0.02396436, -0.2993668, 0.018079046, 0.0123179965, 0.019356515, -0.3041985, 0.0026812062, 0.005565926, 0.015305976, -0.30212662, -0.009646894, 7.446508e-05, 0.011778627, -0.2945912, -0.019287577, -0.0043050377, 0.00873708, -0.28284675, -0.026597979, -0.007712748, 0.00614207}};
	localparam real hf[0:1199] = {0.08329454, -0.002166092, -0.0027761427, 0.00011518025, 0.08110477, -0.0063688783, -0.0024798503, 0.00033087053, 0.07689949, -0.010223132, -0.0019210777, 0.0005066809, 0.07090005, -0.013547321, -0.0011514168, 0.00062490307, 0.063409075, -0.016198227, -0.0002336508, 0.0006753596, 0.054789472, -0.018077407, 0.0007636957, 0.00065492233, 0.045441262, -0.019134235, 0.0017715159, 0.00056670024, 0.0357776, -0.0193657, 0.0027247295, 0.00041897726, 0.026201675, -0.01881328, 0.0035661354, 0.00022398416, 0.017085839, -0.017557386, 0.004249371, -3.4112024e-06, 0.008753973, -0.015709942, 0.0047409004, -0.0002470124, 0.0014679186, -0.013405709, 0.0050210143, -0.0004905292, -0.0045815906, -0.010792999, 0.005083893, -0.00071867666, -0.009279324, -0.008024375, 0.0049368176, -0.0009180901, -0.012585424, -0.005247892, 0.004598668, -0.0010780233, -0.014531144, -0.0025993309, 0.0040978594, -0.0011908124, -0.015211031, -0.00019580046, 0.003469903, -0.0012521034, -0.014772323, 0.0018690547, 0.0027547646, -0.0012608538, -0.013402386, 0.003528106, 0.001994197, -0.0012191334, -0.011315072, 0.0047420333, 0.0012292054, -0.0011317527, -0.008736865, 0.0054989457, 0.0004977813, -0.0010057626, -0.0058936058, 0.0058124997, -0.0001669889, -0.0008498637, -0.0029984799, 0.0057187625, -0.000738365, -0.0006737709, -0.00024183313, 0.0052721114, -0.0011969025, -0.00048757452, 0.0022167892, 0.00454049, -0.0015309008, -0.0003011352, 0.0042541414, 0.0036003485, -0.0017363714, -0.00012354564, 0.005786239, 0.0025315832, -0.0018165703, 3.731639e-05, 0.006768852, 0.0014127643, -0.0017811633, 0.0001751257, 0.007195743, 0.0003168895, -0.0016451057, 0.00028532883, 0.0070949555, -0.0006921433, -0.0014273255, 0.00036524286, 0.0065235584, -0.0015622124, -0.0011493044, 0.00041403915, 0.0055612777, -0.0022547294, -0.0008336459, 0.0004326236, 0.0043034963, -0.0027454633, -0.0005027143, 0.00042342985, 0.0028540604, -0.0030244729, -0.000177414, 0.00039014494, 0.0013183362, -0.0030952408, 0.00012383409, 0.00033738976, -0.0002031292, -0.0029731286, 0.00038587966, 0.00027037621, -0.0016200356, -0.0026833103, 0.00059737125, 0.00019456302, -0.002856627, -0.0022583492, 0.0007510202, 0.00011532953, -0.003854726, -0.0017355902, 0.00084361015, 3.76848e-05, -0.0045754556, -0.001154535, 0.0008757757, -3.3975284e-05, -0.0049996753, -0.0005543484, 0.00085158495, -9.6053416e-05, -0.005127238, 2.837238e-05, 0.0007779675, -0.00014587368, -0.004975216, 0.00056146574, 0.0006640366, -0.00018174076, -0.0045753065, 0.0010186381, 0.0005203518, -0.00020293827, -0.0039706375, 0.0013804217, 0.00035817196, -0.00020967193, -0.0032122214, 0.0016346483, 0.00018874014, -0.00020296614, -0.0023552885, 0.0017764589, 2.263921e-05, -0.00018452431, -0.0014557238, 0.0018078935, -0.00013075274, -0.00015656414, -0.00056680525, 0.0017371231, -0.00026368542, -0.00012163978, 0.0002636046, 0.0015774048, -0.0003703254, -8.2462095e-05, 0.0009952903, 0.0013458435, -0.0004469077, -4.1727493e-05, 0.0015972689, 0.0010620521, -0.00049175444, -1.964157e-06, 0.0020486964, 0.0007467939, -0.00050517224, 3.459715e-05, 0.0023391126, 0.00042068918, -0.00048924563, 6.612282e-05, 0.0024680665, 0.000103051025, -0.0004475487, 9.124376e-05, 0.002444209, -0.00018909262, -0.0003847991, 0.000109089655, 0.0022839506, -0.00044175467, -0.0003064791, 0.0001192914, 0.0020098023, -0.0006444992, -0.00021844968, 0.00012195457, 0.0016485278, -0.0007907008, -0.00012657914, 0.000117608244, 0.001229226, -0.00087756186, -3.6406847e-05, 0.00010713449, 0.00078146264, -0.00090591045, 4.7142166e-05, 9.168434e-05, 0.00033355152, -0.00087981, 0.00011998062, 7.2586394e-05, -8.893034e-05, -0.00080602197, 0.00017901315, 5.1253974e-05, -0.00046433104, -0.0006933657, 0.00022221931, 2.9096242e-05, -0.0007757765, -0.00055202167, 0.00024866723, 7.438023e-06, -0.0010116705, -0.0003928233, 0.0002584639, -1.2547952e-05, -0.0011658471, -0.00022657894, 0.00025265085, -2.9893668e-05, -0.0012373996, -6.345961e-05, 0.00023305652, -4.3871765e-05, -0.0012302273, 8.751874e-05, 0.00020211759, -5.401432e-05, -0.0011523513, 0.00021889791, 0.0001626827, -6.011504e-05, -0.0010150615, 0.00032505317, 0.0001178113, -6.2216306e-05, -0.00083195925, 0.0004023383, 7.05795e-05, -6.0583283e-05, -0.0006179596, 0.00044910403, 2.3903529e-05, -5.566773e-05, -0.000388314, 0.00046560107, -1.9611043e-05, -4.8064652e-05, -0.00015770759, 0.00045378428, -5.7787965e-05, -3.8464852e-05, 6.0525042e-05, 0.00041703798, -8.896328e-05, -2.7606573e-05, 0.00025503212, 0.00035984657, -0.00011203119, -1.6228969e-05, 0.00041690344, 0.00028743348, -0.00012645379, -5.0299927e-06, 0.00053994585, 0.00020539254, -0.00013223746, 5.3693966e-06, 0.00062077766, 0.000119333505, -0.00012988062, 1.4453233e-05, 0.0006587534, 3.456041e-05, -0.00012029824, 2.1829897e-05, 0.0006557397, -4.4201966e-05, -0.00010473003, 2.7242548e-05, 0.00061576907, -0.00011302245, -8.463867e-05, 3.057088e-05, 0.00054460356, -0.00016891213, -6.160515e-05, 3.1824948e-05, 0.0004492405, -0.00020990512, -3.7227335e-05, 3.113213e-05, 0.00033739573, -0.00023507322, -1.3027222e-05, 2.8718683e-05, 0.00021699451, -0.00024448003, 9.628657e-06, 2.4887378e-05, 9.569915e-05, -0.00023908276, 2.9592326e-05, 1.999295e-05, -1.9503277e-05, -0.00022059261, 4.5979014e-05, 1.4416896e-05, -0.00012263555, -0.00019130523, 5.8192527e-05, 8.543174e-06, -0.00020897533, -0.00015391411, 6.5931745e-05, 2.736059e-06, -0.00027520536, -0.00011131903, 6.9179645e-05, -2.6787536e-06, -0.00031946908, -6.644102e-05, 6.817724e-05, -7.429047e-06, -0.00034133776, -2.2053635e-05, 6.338518e-05, -1.1306511e-05, -0.0003416992, 1.9361161e-05, 5.543659e-05, -1.41725295e-05, -0.00032258194, 5.572686e-05, 4.508447e-05, -1.5959447e-05, -0.00028693117, 8.545225e-05, 3.3147346e-05, -1.666766e-05, -0.00023835365, 0.00010747597, 2.0456324e-05, -1.6359112e-05, -0.00018084924, 0.00012127665, 7.8064695e-06, -1.51478835e-05, -0.00011854544, 0.00012685123, -4.0851087e-06, -1.3188726e-05, -5.5450007e-05, 0.00012466582, -1.46127495e-05, -1.0664356e-05, 4.7660674e-06, 0.00011558446, -2.3306176e-05, -7.772356e-06, 5.8945756e-05, 0.00010078198, -2.9844436e-05, -4.712502e-06, 0.000104577, 8.164745e-05, -3.4059987e-05, -1.6751434e-06, 0.00013987445, 5.9684568e-05, -3.593366e-05, 1.1687506e-06, 0.00016381207, 3.641501e-05, -3.5581612e-05, 3.6755025e-06, 0.00017610924, 1.32899795e-05, -3.323585e-05, 5.734323e-06, 0.00017717574, -8.385832e-06, -2.9219946e-05, 7.270502e-06, 0.00016802263, -2.7514678e-05, -2.3921879e-05, 8.246232e-06, 0.00015014727, -4.3248623e-05, -1.7765786e-05, 8.659256e-06, 0.00012540168, -5.5014116e-05, -1.1184327e-05, 8.5396105e-06, 9.5853036e-05, -6.2518535e-05, -4.593211e-06, 7.944839e-06, 6.3645406e-05, -6.574011e-05, 1.6309002e-06, 6.954094e-06, 3.0870076e-05, -6.4903375e-05, 7.168145e-06, 5.6615645e-06, -5.486277e-07, -6.0442904e-05, 1.1768293e-05, 4.169675e-06, -2.894718e-05, -5.2958494e-05, 1.5258382e-05, 2.5824618e-06, -5.2992873e-05, -4.3165244e-05, 1.7545217e-05, 9.994867e-07, -7.172828e-05, -3.1841784e-05, 1.8613091e-05, -4.894133e-07, -8.459013e-05, -1.9779827e-05, 1.8517301e-05, -1.8083222e-06, -9.140385e-05, -7.737765e-06, 1.7374226e-05, -2.8982477e-06, -9.235647e-05, 3.5993999e-06, 1.5348875e-05, -3.7188734e-06, -8.795159e-05, 1.3652127e-05, 1.2640844e-05, -4.2490783e-06, -7.895036e-05, 2.1969343e-05, 9.469648e-06, -4.486313e-06, -6.630368e-05, 2.8241926e-05, 6.0602943e-06, -4.444977e-06, -5.107978e-05, 3.2306812e-05, 2.6299333e-06, -4.153981e-06, -3.439219e-05, 3.4142384e-05, -6.2377325e-07, -3.6537178e-06, -1.7331871e-05, 3.3856228e-05, -3.5320716e-06, -2.9926648e-06, -9.0717117e-07, 3.1666685e-05, -5.9619833e-06, -2.2238494e-06, 1.4005824e-05, 2.787986e-05, -7.820482e-06, -1.4013922e-06, 2.6700658e-05, 2.28638e-05, -9.055991e-06, -5.773156e-07, 3.666464e-05, 1.7021604e-05, -9.657375e-06, 2.0122168e-07, 4.358963e-05, 1.0765095e-05, -9.650729e-06, 8.941513e-07, 4.7370126e-05, 4.490504e-06, -9.094336e-06, 1.4701044e-06, 4.808999e-05, -1.4426392e-06, -8.072279e-06, 1.9073723e-06, 4.5999634e-05, -6.7285173e-06, -6.6871944e-06, 2.194223e-06, 4.1485862e-05, -1.1127348e-05, -5.052642e-06, 2.3286218e-06, 3.5036843e-05, -1.4472771e-05, -3.2855949e-06, 2.3174214e-06, 2.7204609e-05, -1.667434e-05, -1.4994419e-06, 2.1751262e-06, 1.8567493e-05, -1.771545e-05, 2.021381e-07, 1.9223355e-06, 9.694645e-06, -1.7647259e-05, 1.7301634e-06, 1.5839881e-06, 1.1144524e-06, -1.6579304e-05, 3.0140243e-06, 1.1875272e-06, -6.7117116e-06, -1.4667707e-05, 4.0037603e-06, 7.6109626e-07, -1.3409413e-05, -1.2101825e-05, 4.6709415e-06, 3.3186762e-07, -1.8704233e-05, -9.090292e-06, 5.008241e-06, -7.541465e-08, -2.2427885e-05, -5.8472865e-06, 5.0278404e-06, -4.396146e-07, -2.4517707e-05, -2.5797851e-06, 4.7588796e-06, -7.440662e-07, -2.5010173e-05, 5.2355216e-07, 4.2441784e-06, -9.770978e-07, -2.4029374e-05, 3.3013955e-06, 3.5364915e-06, -1.1322225e-06, -2.1771586e-05, 5.6263434e-06, 2.6945547e-06, -1.2080135e-06, -1.8487219e-05, 7.4089544e-06, 1.7791652e-06, -1.2077045e-06, -1.4461363e-05, 8.599235e-06, 8.4951876e-07, -1.1385607e-06, -9.994244e-06, 9.18573e-06, -4.0014346e-08, -1.0110807e-06, -5.3826448e-06, 9.192508e-06, -8.4252963e-07, -8.3809e-07, -9.0332435e-07, 8.674402e-06, -1.5205522e-06, -6.337877e-07, 3.2008677e-06, 7.710956e-06, -2.047276e-06, -4.128062e-07, 6.731606e-06, 6.3995335e-06, -2.4070757e-06, -1.8933547e-07, 9.542158e-06, 4.8480665e-06, -2.5953334e-06, 2.36442e-08, 1.154084e-05, 3.1678962e-06, -2.6176535e-06, 2.1498701e-07, 1.2690999e-05, 1.4670982e-06, -2.4885692e-06, 3.7584263e-07, 1.30078615e-05, -1.5537056e-07, -2.2298634e-06, 4.9994225e-07, 1.2552728e-05, -1.614445e-06, -1.8686356e-06, 5.837101e-07, 1.1425081e-05, -2.8424806e-06, -1.4352513e-06, 6.2621103e-07, 9.753283e-06, -3.7914517e-06, -9.61298e-07, 6.289522e-07, 7.6845e-06, -4.433821e-06, -4.7766804e-07, 5.955645e-07, 5.3745202e-06, -4.762158e-06, -1.2863228e-08, 5.3139325e-07, 2.9780485e-06, -4.78765e-06, 4.0840303e-07, 4.430303e-07, 6.3998715e-07, -4.537688e-06, 7.6625406e-07, 3.378189e-07, -1.5118944e-06, -4.0527616e-06, 1.046323e-06, 2.2336387e-07, -3.372613e-06, -3.3829053e-06, 1.2400466e-06, 1.0707267e-07, -4.8637894e-06, -2.5839322e-06, 1.3446019e-06, -4.248001e-09, -5.935583e-06, -1.7137032e-06, 1.3625194e-06, -1.04723284e-07, -6.566817e-06, -8.2863176e-07, 1.3010292e-06, -1.8965635e-07, -6.7634546e-06, 1.939584e-08, 1.1712015e-06, -2.5568409e-07, -6.555675e-06, 7.855475e-07, 9.869489e-07, -3.008418e-07, -5.993846e-06, 1.4339305e-06, 7.639624e-07, -3.245421e-07, -5.143728e-06, 1.9387867e-06, 5.186478e-07, -3.274772e-07, -4.0812574e-06, 2.284996e-06, 2.671212e-07, -3.1145754e-07, -2.8872491e-06, 2.4679262e-06, 2.431808e-08, -2.7920208e-07, -1.6423209e-06, 2.4926965e-06, -1.9674613e-07, -2.3409666e-07, -4.2231613e-07, 2.372959e-06, -3.8553537e-07, -1.7993743e-07, 7.0556695e-07, 2.1293054e-06, -5.343577e-07, -1.2067527e-07, 1.6857839e-06, 1.7874331e-06, -6.385329e-07, -6.017576e-08, 2.4765015e-06, 1.3761929e-06, -6.963727e-07, -2.0068598e-09, 3.0506776e-06, 9.2564335e-07, -7.08992e-07, 5.0736222e-08, 3.3961942e-06, 4.6522177e-07, -6.7997814e-07, 9.55625e-08, 3.515127e-06, 2.212465e-08, -6.1495115e-07, 1.3066972e-07, 3.4222758e-06, -3.800299e-07, -5.210494e-07, 1.5498154e-07, 3.1431073e-06, -7.222081e-07, -4.0637804e-07, 1.6813975e-07, 2.711288e-06, -9.906094e-07, -2.7945455e-07, 1.7045632e-07, 2.165983e-06, -1.1769547e-06, -1.4868394e-07, 1.6283175e-07, 1.5490983e-06, -1.2784332e-06, -2.1890017e-08, 1.4664774e-07, 9.026308e-07, -1.2973412e-06, 9.407538e-08, 1.2364242e-07, 2.6626404e-07, -1.2404652e-06, 1.9363054e-07, 9.5777445e-08, -3.2467412e-07, -1.1182668e-06, 2.7266123e-07, 6.510469e-08, -8.408114e-07, -9.439365e-07, 3.2861544e-07, 3.3640767e-08, -1.2598389e-06, -7.323812e-07, 3.6050037e-07, 3.2552991e-09, -1.5671101e-06, -4.9921067e-07, 3.6879018e-07, -2.4421656e-08, -1.7557471e-06, -2.5978076e-07, 3.5525957e-07, -4.8069758e-08, -1.8262921e-06, -2.834151e-08, 3.2275847e-07, -6.6724176e-08, -1.78597e-06, 1.8266994e-07, 2.7494718e-07, -7.979675e-08, -1.6476401e-06, 3.6316598e-07, 2.1601049e-07, -8.707365e-08, -1.4285262e-06, 5.0576006e-07, 1.5036903e-07, -8.869193e-08, -1.1488177e-06, 6.0593055e-07, 8.240474e-08, -8.5098264e-08, -8.302372e-07, 6.6200585e-07, 1.621461e-08, -7.699403e-08, -4.946546e-07, 6.749881e-07, -4.4595726e-08, -6.527098e-08, -1.628267e-07, 6.482414e-07, -9.7070874e-08, -5.094235e-08, 1.4668123e-07, 5.8707514e-07, -1.3901226e-07, -3.5073416e-08, 4.183448e-07, 4.982559e-07, -1.6903141e-07, -1.8715838e-08, 6.4027654e-07, 3.8948244e-07, -1.86552e-07, -2.848981e-09, 8.0455715e-07, 2.6885849e-07, -1.9176534e-07, 1.1669062e-08, 9.073094e-07, 1.4439148e-07, -1.8554638e-07, 2.4138847e-08, 9.485341e-07, 2.3545416e-08, -1.6933865e-07, 3.4044355e-08, 9.317406e-07, -8.713313e-08, -1.4501784e-07, 4.106495e-08, 8.6341265e-07, -1.8230097e-07, -1.1474362e-07, 4.507505e-08, 7.523552e-07, -2.5800833e-07, -8.0809485e-08, 4.6132715e-08, 6.089715e-07, -3.1179144e-07, -4.5499178e-08, 4.445884e-08, 4.4451713e-07, -3.4267146e-07, -1.0957408e-08, 4.0409056e-08, 2.7037726e-07, -3.5106885e-07, 2.091922e-08, 3.4440603e-08, 9.7405064e-08, -3.3864612e-07, 4.856674e-08, 2.7076597e-08, -6.464668e-08, -3.080948e-07, 7.081131e-08, 1.8869901e-08, -2.0757685e-07, -2.6288382e-07, 8.689902e-08, 1.03687805e-08, -3.2505588e-07, -2.0698765e-07, 9.6498866e-08, 2.0860698e-09, -4.1280853e-07, -1.4461165e-07, 9.9681344e-08, -5.5266987e-09, -4.6866188e-07, -7.993008e-08, 9.687621e-08, -1.2099203e-08, -4.9246916e-07, -1.6851118e-08, 8.881373e-08, -1.7355719e-08, -4.8592494e-07, 4.118071e-08, 7.645443e-08, -2.112183e-08, -4.5229345e-07, 9.133676e-08, 6.0912384e-08, -2.332472e-08, -3.9607247e-07, 1.3150695e-07, 4.3377042e-08, -2.3987662e-08, -3.226197e-07, 1.6035165e-07, 2.503825e-08, -2.3219524e-08, -2.3776522e-07, 1.7730463e-07, 7.018331e-09, -2.120042e-08, -1.4743395e-07, 1.825318e-07, -9.685473e-09, -1.816464e-08, -5.7298827e-08, 1.7685193e-07, -2.4245953e-08, -1.4382141e-08, 2.751871e-08, 1.6162778e-07, -3.6036923e-08, -1.013975e-08, 1.026883e-07, 1.386366e-07, -4.464977e-08, -5.7231997e-09, 1.648422e-07, 1.09929275e-07, -4.989604e-08, -1.4009387e-09, 2.1167571e-07, 7.768735e-08, -5.1797212e-08, 2.5895295e-09, 2.419773e-07, 4.4086146e-08, -5.0563482e-08, 6.052244e-09, 2.5559356e-07, 1.1171274e-08, -4.6563798e-08, 8.840005e-09, 2.5333728e-07, -1.9245604e-08, -4.028969e-08, 1.0858124e-08, 2.368489e-07, -4.5667843e-08, -3.2315594e-08, 1.206482e-08, 2.084243e-07, -6.696915e-08, -2.3258158e-08, 1.2468566e-08, 1.7082131e-07, -8.242253e-08, -1.3737084e-08, 1.2122815e-08, 1.2705854e-07, -9.170374e-08, -4.3394865e-09, 1.1118672e-08, 8.0218335e-08, -9.487138e-08, 4.410481e-09, 9.5761115e-09, 3.3264943e-08, -9.232712e-08, 1.2075523e-08, 7.634381e-09, -1.1113255e-08, -8.476008e-08, 1.8321863e-08, 5.442233e-09, -5.06308e-08, -7.3080194e-08, 2.292842e-08, 3.1485288e-09, -8.34971e-08, -5.8345268e-08, 2.5788685e-08, 8.937436e-10, -1.0847142e-07, -4.168657e-08, 2.6905875e-08, -1.1972464e-09, -1.2488124e-07, -2.4237318e-08, 2.6382303e-08, -3.0208003e-09, -1.326065e-07, -7.067889e-09, 2.4404104e-08, -4.4983994e-09, -1.3203386e-07, 8.869257e-09, 2.122264e-08, -5.578732e-09, -1.239863e-07, 2.2782649e-08, 1.7133946e-08, -6.23803e-09, -1.0963473e-07, 3.407161e-08, 1.2457596e-08, -6.478797e-09, -9.039801e-08, 4.234234e-08, 7.516241e-09, -6.3271677e-09, -6.7838435e-08, 4.741066e-08, 2.6169107e-09, -5.8291634e-09, -4.3559e-08, 4.9292566e-08, -1.965005e-09, -5.046175e-09, -1.9108095e-08, 4.8184237e-08, -5.9984484e-09, -4.0499977e-09, 4.1036015e-09, 4.4433687e-08, -9.305645e-09, -2.9177456e-09, 2.4870431e-08, 3.850646e-08, -1.1767171e-08, -1.7269481e-09, 4.2241e-08, 3.0947895e-08, -1.3323201e-08, -5.510889e-10, 5.5548206e-08, 2.2344404e-08, -1.39712455e-08, 5.441997e-10, 6.4420206e-08, 1.3286148e-08, -1.3760832e-08, 1.5041312e-09, 6.877351e-08, 4.333001e-09, -1.2785725e-08, 2.2868563e-09, 6.879024e-08, -4.014479e-09, -1.1174368e-08, 2.864617e-09, 6.488251e-08, -1.1337952e-08, -9.079252e-09, 3.2239882e-09, 5.7646943e-08, -1.731732e-08, -6.66593e-09, 3.3652767e-09, 4.7813135e-08, -2.1739618e-08, -4.102335e-09, 3.3011978e-09, 3.6189345e-08, -2.4500967e-08, -1.5489727e-09, 3.0549656e-09, 2.3608933e-08, -2.5602098e-08, 8.495212e-10, 2.657972e-09, 1.0880434e-08, -2.5138347e-08, 2.9711198e-09, 2.147216e-09, -1.2561846e-09, -2.328521e-08, 4.7212088e-09, 1.5626592e-09, -1.2165187e-08, -2.0280703e-08, 6.0353718e-09, 9.446669e-10, -2.1341396e-08, -1.6405826e-08, 6.880187e-09, 3.3166533e-10, -2.8426568e-08, -1.1964452e-08, 7.252182e-09, -2.418632e-10, -3.3215823e-08, -7.263813e-09, 7.175178e-09, -7.4697204e-10, -3.565473e-08, -2.5966669e-09, 6.696332e-09, -1.1613733e-09, -3.5828066e-08, 1.7740251e-09, 5.8812253e-09, -1.4700747e-09, -3.3941735e-08, 5.6272538e-09, 4.8083684e-09, -1.6655398e-09, -3.0299493e-08, 8.792569e-09, 3.5634935e-09, -1.7474071e-09, -2.5276282e-08, 1.1154986e-08, 2.2339752e-09, -1.721828e-09, -1.9290098e-08, 1.2656258e-08, 9.0369406e-10, -1.6004952e-09, -1.2774032e-08, 1.32927935e-08, -3.5141617e-10, -1.3994481e-09, -6.1501435e-09, 1.31106574e-08, -1.4669405e-09, -1.1377443e-09, 1.9355972e-10, 1.2198212e-08, -2.3925593e-09, -8.360854e-10, 5.922004e-09, 1.0677051e-08, -3.0935758e-09, -5.154796e-10, 1.0767118e-08, 8.6919005e-09, -3.551406e-09, -1.9601447e-10, 1.45367345e-08, 6.40016e-09, -3.7631045e-09, 1.0420049e-10, 1.7118325e-08, 3.961722e-09, -3.740042e-09, 3.6987857e-10, 1.8477824e-08, 1.5296149e-09, -3.505894e-09, 5.891586e-10, 1.8654106e-08, -7.5806944e-10, -3.0941185e-09, 7.5395507e-10, 1.7749816e-08, -2.7846279e-09, -2.5451163e-09, 8.600596e-10, 1.5919445e-08, -4.459364e-09, -1.9032655e-09, 9.070116e-10, 1.335558e-08, -5.7202834e-09, -1.2140127e-09, 8.977677e-10, 1.0274292e-08, -6.5348953e-09, -5.2117805e-10, 8.3820756e-10, 6.9005788e-09, -6.899254e-09, 1.3538694e-10, 7.3652023e-10, 3.4546863e-09, -6.8354673e-09, 7.216952e-10, 6.0251704e-10, 1.3999661e-10, -6.3879524e-09, 1.2110034e-09, 4.4691778e-10, -2.8669613e-09, -5.6187783e-09, 1.5846467e-09, 2.806527e-10, -5.4240217e-09, -4.602446e-09, 1.8323345e-09, 1.1421921e-10};
	localparam real hb[0:1199] = {0.08329454, 0.002166092, -0.0027761427, -0.00011518025, 0.08110477, 0.0063688783, -0.0024798503, -0.00033087053, 0.07689949, 0.010223132, -0.0019210777, -0.0005066809, 0.07090005, 0.013547321, -0.0011514168, -0.00062490307, 0.063409075, 0.016198227, -0.0002336508, -0.0006753596, 0.054789472, 0.018077407, 0.0007636957, -0.00065492233, 0.045441262, 0.019134235, 0.0017715159, -0.00056670024, 0.0357776, 0.0193657, 0.0027247295, -0.00041897726, 0.026201675, 0.01881328, 0.0035661354, -0.00022398416, 0.017085839, 0.017557386, 0.004249371, 3.4112024e-06, 0.008753973, 0.015709942, 0.0047409004, 0.0002470124, 0.0014679186, 0.013405709, 0.0050210143, 0.0004905292, -0.0045815906, 0.010792999, 0.005083893, 0.00071867666, -0.009279324, 0.008024375, 0.0049368176, 0.0009180901, -0.012585424, 0.005247892, 0.004598668, 0.0010780233, -0.014531144, 0.0025993309, 0.0040978594, 0.0011908124, -0.015211031, 0.00019580046, 0.003469903, 0.0012521034, -0.014772323, -0.0018690547, 0.0027547646, 0.0012608538, -0.013402386, -0.003528106, 0.001994197, 0.0012191334, -0.011315072, -0.0047420333, 0.0012292054, 0.0011317527, -0.008736865, -0.0054989457, 0.0004977813, 0.0010057626, -0.0058936058, -0.0058124997, -0.0001669889, 0.0008498637, -0.0029984799, -0.0057187625, -0.000738365, 0.0006737709, -0.00024183313, -0.0052721114, -0.0011969025, 0.00048757452, 0.0022167892, -0.00454049, -0.0015309008, 0.0003011352, 0.0042541414, -0.0036003485, -0.0017363714, 0.00012354564, 0.005786239, -0.0025315832, -0.0018165703, -3.731639e-05, 0.006768852, -0.0014127643, -0.0017811633, -0.0001751257, 0.007195743, -0.0003168895, -0.0016451057, -0.00028532883, 0.0070949555, 0.0006921433, -0.0014273255, -0.00036524286, 0.0065235584, 0.0015622124, -0.0011493044, -0.00041403915, 0.0055612777, 0.0022547294, -0.0008336459, -0.0004326236, 0.0043034963, 0.0027454633, -0.0005027143, -0.00042342985, 0.0028540604, 0.0030244729, -0.000177414, -0.00039014494, 0.0013183362, 0.0030952408, 0.00012383409, -0.00033738976, -0.0002031292, 0.0029731286, 0.00038587966, -0.00027037621, -0.0016200356, 0.0026833103, 0.00059737125, -0.00019456302, -0.002856627, 0.0022583492, 0.0007510202, -0.00011532953, -0.003854726, 0.0017355902, 0.00084361015, -3.76848e-05, -0.0045754556, 0.001154535, 0.0008757757, 3.3975284e-05, -0.0049996753, 0.0005543484, 0.00085158495, 9.6053416e-05, -0.005127238, -2.837238e-05, 0.0007779675, 0.00014587368, -0.004975216, -0.00056146574, 0.0006640366, 0.00018174076, -0.0045753065, -0.0010186381, 0.0005203518, 0.00020293827, -0.0039706375, -0.0013804217, 0.00035817196, 0.00020967193, -0.0032122214, -0.0016346483, 0.00018874014, 0.00020296614, -0.0023552885, -0.0017764589, 2.263921e-05, 0.00018452431, -0.0014557238, -0.0018078935, -0.00013075274, 0.00015656414, -0.00056680525, -0.0017371231, -0.00026368542, 0.00012163978, 0.0002636046, -0.0015774048, -0.0003703254, 8.2462095e-05, 0.0009952903, -0.0013458435, -0.0004469077, 4.1727493e-05, 0.0015972689, -0.0010620521, -0.00049175444, 1.964157e-06, 0.0020486964, -0.0007467939, -0.00050517224, -3.459715e-05, 0.0023391126, -0.00042068918, -0.00048924563, -6.612282e-05, 0.0024680665, -0.000103051025, -0.0004475487, -9.124376e-05, 0.002444209, 0.00018909262, -0.0003847991, -0.000109089655, 0.0022839506, 0.00044175467, -0.0003064791, -0.0001192914, 0.0020098023, 0.0006444992, -0.00021844968, -0.00012195457, 0.0016485278, 0.0007907008, -0.00012657914, -0.000117608244, 0.001229226, 0.00087756186, -3.6406847e-05, -0.00010713449, 0.00078146264, 0.00090591045, 4.7142166e-05, -9.168434e-05, 0.00033355152, 0.00087981, 0.00011998062, -7.2586394e-05, -8.893034e-05, 0.00080602197, 0.00017901315, -5.1253974e-05, -0.00046433104, 0.0006933657, 0.00022221931, -2.9096242e-05, -0.0007757765, 0.00055202167, 0.00024866723, -7.438023e-06, -0.0010116705, 0.0003928233, 0.0002584639, 1.2547952e-05, -0.0011658471, 0.00022657894, 0.00025265085, 2.9893668e-05, -0.0012373996, 6.345961e-05, 0.00023305652, 4.3871765e-05, -0.0012302273, -8.751874e-05, 0.00020211759, 5.401432e-05, -0.0011523513, -0.00021889791, 0.0001626827, 6.011504e-05, -0.0010150615, -0.00032505317, 0.0001178113, 6.2216306e-05, -0.00083195925, -0.0004023383, 7.05795e-05, 6.0583283e-05, -0.0006179596, -0.00044910403, 2.3903529e-05, 5.566773e-05, -0.000388314, -0.00046560107, -1.9611043e-05, 4.8064652e-05, -0.00015770759, -0.00045378428, -5.7787965e-05, 3.8464852e-05, 6.0525042e-05, -0.00041703798, -8.896328e-05, 2.7606573e-05, 0.00025503212, -0.00035984657, -0.00011203119, 1.6228969e-05, 0.00041690344, -0.00028743348, -0.00012645379, 5.0299927e-06, 0.00053994585, -0.00020539254, -0.00013223746, -5.3693966e-06, 0.00062077766, -0.000119333505, -0.00012988062, -1.4453233e-05, 0.0006587534, -3.456041e-05, -0.00012029824, -2.1829897e-05, 0.0006557397, 4.4201966e-05, -0.00010473003, -2.7242548e-05, 0.00061576907, 0.00011302245, -8.463867e-05, -3.057088e-05, 0.00054460356, 0.00016891213, -6.160515e-05, -3.1824948e-05, 0.0004492405, 0.00020990512, -3.7227335e-05, -3.113213e-05, 0.00033739573, 0.00023507322, -1.3027222e-05, -2.8718683e-05, 0.00021699451, 0.00024448003, 9.628657e-06, -2.4887378e-05, 9.569915e-05, 0.00023908276, 2.9592326e-05, -1.999295e-05, -1.9503277e-05, 0.00022059261, 4.5979014e-05, -1.4416896e-05, -0.00012263555, 0.00019130523, 5.8192527e-05, -8.543174e-06, -0.00020897533, 0.00015391411, 6.5931745e-05, -2.736059e-06, -0.00027520536, 0.00011131903, 6.9179645e-05, 2.6787536e-06, -0.00031946908, 6.644102e-05, 6.817724e-05, 7.429047e-06, -0.00034133776, 2.2053635e-05, 6.338518e-05, 1.1306511e-05, -0.0003416992, -1.9361161e-05, 5.543659e-05, 1.41725295e-05, -0.00032258194, -5.572686e-05, 4.508447e-05, 1.5959447e-05, -0.00028693117, -8.545225e-05, 3.3147346e-05, 1.666766e-05, -0.00023835365, -0.00010747597, 2.0456324e-05, 1.6359112e-05, -0.00018084924, -0.00012127665, 7.8064695e-06, 1.51478835e-05, -0.00011854544, -0.00012685123, -4.0851087e-06, 1.3188726e-05, -5.5450007e-05, -0.00012466582, -1.46127495e-05, 1.0664356e-05, 4.7660674e-06, -0.00011558446, -2.3306176e-05, 7.772356e-06, 5.8945756e-05, -0.00010078198, -2.9844436e-05, 4.712502e-06, 0.000104577, -8.164745e-05, -3.4059987e-05, 1.6751434e-06, 0.00013987445, -5.9684568e-05, -3.593366e-05, -1.1687506e-06, 0.00016381207, -3.641501e-05, -3.5581612e-05, -3.6755025e-06, 0.00017610924, -1.32899795e-05, -3.323585e-05, -5.734323e-06, 0.00017717574, 8.385832e-06, -2.9219946e-05, -7.270502e-06, 0.00016802263, 2.7514678e-05, -2.3921879e-05, -8.246232e-06, 0.00015014727, 4.3248623e-05, -1.7765786e-05, -8.659256e-06, 0.00012540168, 5.5014116e-05, -1.1184327e-05, -8.5396105e-06, 9.5853036e-05, 6.2518535e-05, -4.593211e-06, -7.944839e-06, 6.3645406e-05, 6.574011e-05, 1.6309002e-06, -6.954094e-06, 3.0870076e-05, 6.4903375e-05, 7.168145e-06, -5.6615645e-06, -5.486277e-07, 6.0442904e-05, 1.1768293e-05, -4.169675e-06, -2.894718e-05, 5.2958494e-05, 1.5258382e-05, -2.5824618e-06, -5.2992873e-05, 4.3165244e-05, 1.7545217e-05, -9.994867e-07, -7.172828e-05, 3.1841784e-05, 1.8613091e-05, 4.894133e-07, -8.459013e-05, 1.9779827e-05, 1.8517301e-05, 1.8083222e-06, -9.140385e-05, 7.737765e-06, 1.7374226e-05, 2.8982477e-06, -9.235647e-05, -3.5993999e-06, 1.5348875e-05, 3.7188734e-06, -8.795159e-05, -1.3652127e-05, 1.2640844e-05, 4.2490783e-06, -7.895036e-05, -2.1969343e-05, 9.469648e-06, 4.486313e-06, -6.630368e-05, -2.8241926e-05, 6.0602943e-06, 4.444977e-06, -5.107978e-05, -3.2306812e-05, 2.6299333e-06, 4.153981e-06, -3.439219e-05, -3.4142384e-05, -6.2377325e-07, 3.6537178e-06, -1.7331871e-05, -3.3856228e-05, -3.5320716e-06, 2.9926648e-06, -9.0717117e-07, -3.1666685e-05, -5.9619833e-06, 2.2238494e-06, 1.4005824e-05, -2.787986e-05, -7.820482e-06, 1.4013922e-06, 2.6700658e-05, -2.28638e-05, -9.055991e-06, 5.773156e-07, 3.666464e-05, -1.7021604e-05, -9.657375e-06, -2.0122168e-07, 4.358963e-05, -1.0765095e-05, -9.650729e-06, -8.941513e-07, 4.7370126e-05, -4.490504e-06, -9.094336e-06, -1.4701044e-06, 4.808999e-05, 1.4426392e-06, -8.072279e-06, -1.9073723e-06, 4.5999634e-05, 6.7285173e-06, -6.6871944e-06, -2.194223e-06, 4.1485862e-05, 1.1127348e-05, -5.052642e-06, -2.3286218e-06, 3.5036843e-05, 1.4472771e-05, -3.2855949e-06, -2.3174214e-06, 2.7204609e-05, 1.667434e-05, -1.4994419e-06, -2.1751262e-06, 1.8567493e-05, 1.771545e-05, 2.021381e-07, -1.9223355e-06, 9.694645e-06, 1.7647259e-05, 1.7301634e-06, -1.5839881e-06, 1.1144524e-06, 1.6579304e-05, 3.0140243e-06, -1.1875272e-06, -6.7117116e-06, 1.4667707e-05, 4.0037603e-06, -7.6109626e-07, -1.3409413e-05, 1.2101825e-05, 4.6709415e-06, -3.3186762e-07, -1.8704233e-05, 9.090292e-06, 5.008241e-06, 7.541465e-08, -2.2427885e-05, 5.8472865e-06, 5.0278404e-06, 4.396146e-07, -2.4517707e-05, 2.5797851e-06, 4.7588796e-06, 7.440662e-07, -2.5010173e-05, -5.2355216e-07, 4.2441784e-06, 9.770978e-07, -2.4029374e-05, -3.3013955e-06, 3.5364915e-06, 1.1322225e-06, -2.1771586e-05, -5.6263434e-06, 2.6945547e-06, 1.2080135e-06, -1.8487219e-05, -7.4089544e-06, 1.7791652e-06, 1.2077045e-06, -1.4461363e-05, -8.599235e-06, 8.4951876e-07, 1.1385607e-06, -9.994244e-06, -9.18573e-06, -4.0014346e-08, 1.0110807e-06, -5.3826448e-06, -9.192508e-06, -8.4252963e-07, 8.3809e-07, -9.0332435e-07, -8.674402e-06, -1.5205522e-06, 6.337877e-07, 3.2008677e-06, -7.710956e-06, -2.047276e-06, 4.128062e-07, 6.731606e-06, -6.3995335e-06, -2.4070757e-06, 1.8933547e-07, 9.542158e-06, -4.8480665e-06, -2.5953334e-06, -2.36442e-08, 1.154084e-05, -3.1678962e-06, -2.6176535e-06, -2.1498701e-07, 1.2690999e-05, -1.4670982e-06, -2.4885692e-06, -3.7584263e-07, 1.30078615e-05, 1.5537056e-07, -2.2298634e-06, -4.9994225e-07, 1.2552728e-05, 1.614445e-06, -1.8686356e-06, -5.837101e-07, 1.1425081e-05, 2.8424806e-06, -1.4352513e-06, -6.2621103e-07, 9.753283e-06, 3.7914517e-06, -9.61298e-07, -6.289522e-07, 7.6845e-06, 4.433821e-06, -4.7766804e-07, -5.955645e-07, 5.3745202e-06, 4.762158e-06, -1.2863228e-08, -5.3139325e-07, 2.9780485e-06, 4.78765e-06, 4.0840303e-07, -4.430303e-07, 6.3998715e-07, 4.537688e-06, 7.6625406e-07, -3.378189e-07, -1.5118944e-06, 4.0527616e-06, 1.046323e-06, -2.2336387e-07, -3.372613e-06, 3.3829053e-06, 1.2400466e-06, -1.0707267e-07, -4.8637894e-06, 2.5839322e-06, 1.3446019e-06, 4.248001e-09, -5.935583e-06, 1.7137032e-06, 1.3625194e-06, 1.04723284e-07, -6.566817e-06, 8.2863176e-07, 1.3010292e-06, 1.8965635e-07, -6.7634546e-06, -1.939584e-08, 1.1712015e-06, 2.5568409e-07, -6.555675e-06, -7.855475e-07, 9.869489e-07, 3.008418e-07, -5.993846e-06, -1.4339305e-06, 7.639624e-07, 3.245421e-07, -5.143728e-06, -1.9387867e-06, 5.186478e-07, 3.274772e-07, -4.0812574e-06, -2.284996e-06, 2.671212e-07, 3.1145754e-07, -2.8872491e-06, -2.4679262e-06, 2.431808e-08, 2.7920208e-07, -1.6423209e-06, -2.4926965e-06, -1.9674613e-07, 2.3409666e-07, -4.2231613e-07, -2.372959e-06, -3.8553537e-07, 1.7993743e-07, 7.0556695e-07, -2.1293054e-06, -5.343577e-07, 1.2067527e-07, 1.6857839e-06, -1.7874331e-06, -6.385329e-07, 6.017576e-08, 2.4765015e-06, -1.3761929e-06, -6.963727e-07, 2.0068598e-09, 3.0506776e-06, -9.2564335e-07, -7.08992e-07, -5.0736222e-08, 3.3961942e-06, -4.6522177e-07, -6.7997814e-07, -9.55625e-08, 3.515127e-06, -2.212465e-08, -6.1495115e-07, -1.3066972e-07, 3.4222758e-06, 3.800299e-07, -5.210494e-07, -1.5498154e-07, 3.1431073e-06, 7.222081e-07, -4.0637804e-07, -1.6813975e-07, 2.711288e-06, 9.906094e-07, -2.7945455e-07, -1.7045632e-07, 2.165983e-06, 1.1769547e-06, -1.4868394e-07, -1.6283175e-07, 1.5490983e-06, 1.2784332e-06, -2.1890017e-08, -1.4664774e-07, 9.026308e-07, 1.2973412e-06, 9.407538e-08, -1.2364242e-07, 2.6626404e-07, 1.2404652e-06, 1.9363054e-07, -9.5777445e-08, -3.2467412e-07, 1.1182668e-06, 2.7266123e-07, -6.510469e-08, -8.408114e-07, 9.439365e-07, 3.2861544e-07, -3.3640767e-08, -1.2598389e-06, 7.323812e-07, 3.6050037e-07, -3.2552991e-09, -1.5671101e-06, 4.9921067e-07, 3.6879018e-07, 2.4421656e-08, -1.7557471e-06, 2.5978076e-07, 3.5525957e-07, 4.8069758e-08, -1.8262921e-06, 2.834151e-08, 3.2275847e-07, 6.6724176e-08, -1.78597e-06, -1.8266994e-07, 2.7494718e-07, 7.979675e-08, -1.6476401e-06, -3.6316598e-07, 2.1601049e-07, 8.707365e-08, -1.4285262e-06, -5.0576006e-07, 1.5036903e-07, 8.869193e-08, -1.1488177e-06, -6.0593055e-07, 8.240474e-08, 8.5098264e-08, -8.302372e-07, -6.6200585e-07, 1.621461e-08, 7.699403e-08, -4.946546e-07, -6.749881e-07, -4.4595726e-08, 6.527098e-08, -1.628267e-07, -6.482414e-07, -9.7070874e-08, 5.094235e-08, 1.4668123e-07, -5.8707514e-07, -1.3901226e-07, 3.5073416e-08, 4.183448e-07, -4.982559e-07, -1.6903141e-07, 1.8715838e-08, 6.4027654e-07, -3.8948244e-07, -1.86552e-07, 2.848981e-09, 8.0455715e-07, -2.6885849e-07, -1.9176534e-07, -1.1669062e-08, 9.073094e-07, -1.4439148e-07, -1.8554638e-07, -2.4138847e-08, 9.485341e-07, -2.3545416e-08, -1.6933865e-07, -3.4044355e-08, 9.317406e-07, 8.713313e-08, -1.4501784e-07, -4.106495e-08, 8.6341265e-07, 1.8230097e-07, -1.1474362e-07, -4.507505e-08, 7.523552e-07, 2.5800833e-07, -8.0809485e-08, -4.6132715e-08, 6.089715e-07, 3.1179144e-07, -4.5499178e-08, -4.445884e-08, 4.4451713e-07, 3.4267146e-07, -1.0957408e-08, -4.0409056e-08, 2.7037726e-07, 3.5106885e-07, 2.091922e-08, -3.4440603e-08, 9.7405064e-08, 3.3864612e-07, 4.856674e-08, -2.7076597e-08, -6.464668e-08, 3.080948e-07, 7.081131e-08, -1.8869901e-08, -2.0757685e-07, 2.6288382e-07, 8.689902e-08, -1.03687805e-08, -3.2505588e-07, 2.0698765e-07, 9.6498866e-08, -2.0860698e-09, -4.1280853e-07, 1.4461165e-07, 9.9681344e-08, 5.5266987e-09, -4.6866188e-07, 7.993008e-08, 9.687621e-08, 1.2099203e-08, -4.9246916e-07, 1.6851118e-08, 8.881373e-08, 1.7355719e-08, -4.8592494e-07, -4.118071e-08, 7.645443e-08, 2.112183e-08, -4.5229345e-07, -9.133676e-08, 6.0912384e-08, 2.332472e-08, -3.9607247e-07, -1.3150695e-07, 4.3377042e-08, 2.3987662e-08, -3.226197e-07, -1.6035165e-07, 2.503825e-08, 2.3219524e-08, -2.3776522e-07, -1.7730463e-07, 7.018331e-09, 2.120042e-08, -1.4743395e-07, -1.825318e-07, -9.685473e-09, 1.816464e-08, -5.7298827e-08, -1.7685193e-07, -2.4245953e-08, 1.4382141e-08, 2.751871e-08, -1.6162778e-07, -3.6036923e-08, 1.013975e-08, 1.026883e-07, -1.386366e-07, -4.464977e-08, 5.7231997e-09, 1.648422e-07, -1.09929275e-07, -4.989604e-08, 1.4009387e-09, 2.1167571e-07, -7.768735e-08, -5.1797212e-08, -2.5895295e-09, 2.419773e-07, -4.4086146e-08, -5.0563482e-08, -6.052244e-09, 2.5559356e-07, -1.1171274e-08, -4.6563798e-08, -8.840005e-09, 2.5333728e-07, 1.9245604e-08, -4.028969e-08, -1.0858124e-08, 2.368489e-07, 4.5667843e-08, -3.2315594e-08, -1.206482e-08, 2.084243e-07, 6.696915e-08, -2.3258158e-08, -1.2468566e-08, 1.7082131e-07, 8.242253e-08, -1.3737084e-08, -1.2122815e-08, 1.2705854e-07, 9.170374e-08, -4.3394865e-09, -1.1118672e-08, 8.0218335e-08, 9.487138e-08, 4.410481e-09, -9.5761115e-09, 3.3264943e-08, 9.232712e-08, 1.2075523e-08, -7.634381e-09, -1.1113255e-08, 8.476008e-08, 1.8321863e-08, -5.442233e-09, -5.06308e-08, 7.3080194e-08, 2.292842e-08, -3.1485288e-09, -8.34971e-08, 5.8345268e-08, 2.5788685e-08, -8.937436e-10, -1.0847142e-07, 4.168657e-08, 2.6905875e-08, 1.1972464e-09, -1.2488124e-07, 2.4237318e-08, 2.6382303e-08, 3.0208003e-09, -1.326065e-07, 7.067889e-09, 2.4404104e-08, 4.4983994e-09, -1.3203386e-07, -8.869257e-09, 2.122264e-08, 5.578732e-09, -1.239863e-07, -2.2782649e-08, 1.7133946e-08, 6.23803e-09, -1.0963473e-07, -3.407161e-08, 1.2457596e-08, 6.478797e-09, -9.039801e-08, -4.234234e-08, 7.516241e-09, 6.3271677e-09, -6.7838435e-08, -4.741066e-08, 2.6169107e-09, 5.8291634e-09, -4.3559e-08, -4.9292566e-08, -1.965005e-09, 5.046175e-09, -1.9108095e-08, -4.8184237e-08, -5.9984484e-09, 4.0499977e-09, 4.1036015e-09, -4.4433687e-08, -9.305645e-09, 2.9177456e-09, 2.4870431e-08, -3.850646e-08, -1.1767171e-08, 1.7269481e-09, 4.2241e-08, -3.0947895e-08, -1.3323201e-08, 5.510889e-10, 5.5548206e-08, -2.2344404e-08, -1.39712455e-08, -5.441997e-10, 6.4420206e-08, -1.3286148e-08, -1.3760832e-08, -1.5041312e-09, 6.877351e-08, -4.333001e-09, -1.2785725e-08, -2.2868563e-09, 6.879024e-08, 4.014479e-09, -1.1174368e-08, -2.864617e-09, 6.488251e-08, 1.1337952e-08, -9.079252e-09, -3.2239882e-09, 5.7646943e-08, 1.731732e-08, -6.66593e-09, -3.3652767e-09, 4.7813135e-08, 2.1739618e-08, -4.102335e-09, -3.3011978e-09, 3.6189345e-08, 2.4500967e-08, -1.5489727e-09, -3.0549656e-09, 2.3608933e-08, 2.5602098e-08, 8.495212e-10, -2.657972e-09, 1.0880434e-08, 2.5138347e-08, 2.9711198e-09, -2.147216e-09, -1.2561846e-09, 2.328521e-08, 4.7212088e-09, -1.5626592e-09, -1.2165187e-08, 2.0280703e-08, 6.0353718e-09, -9.446669e-10, -2.1341396e-08, 1.6405826e-08, 6.880187e-09, -3.3166533e-10, -2.8426568e-08, 1.1964452e-08, 7.252182e-09, 2.418632e-10, -3.3215823e-08, 7.263813e-09, 7.175178e-09, 7.4697204e-10, -3.565473e-08, 2.5966669e-09, 6.696332e-09, 1.1613733e-09, -3.5828066e-08, -1.7740251e-09, 5.8812253e-09, 1.4700747e-09, -3.3941735e-08, -5.6272538e-09, 4.8083684e-09, 1.6655398e-09, -3.0299493e-08, -8.792569e-09, 3.5634935e-09, 1.7474071e-09, -2.5276282e-08, -1.1154986e-08, 2.2339752e-09, 1.721828e-09, -1.9290098e-08, -1.2656258e-08, 9.0369406e-10, 1.6004952e-09, -1.2774032e-08, -1.32927935e-08, -3.5141617e-10, 1.3994481e-09, -6.1501435e-09, -1.31106574e-08, -1.4669405e-09, 1.1377443e-09, 1.9355972e-10, -1.2198212e-08, -2.3925593e-09, 8.360854e-10, 5.922004e-09, -1.0677051e-08, -3.0935758e-09, 5.154796e-10, 1.0767118e-08, -8.6919005e-09, -3.551406e-09, 1.9601447e-10, 1.45367345e-08, -6.40016e-09, -3.7631045e-09, -1.0420049e-10, 1.7118325e-08, -3.961722e-09, -3.740042e-09, -3.6987857e-10, 1.8477824e-08, -1.5296149e-09, -3.505894e-09, -5.891586e-10, 1.8654106e-08, 7.5806944e-10, -3.0941185e-09, -7.5395507e-10, 1.7749816e-08, 2.7846279e-09, -2.5451163e-09, -8.600596e-10, 1.5919445e-08, 4.459364e-09, -1.9032655e-09, -9.070116e-10, 1.335558e-08, 5.7202834e-09, -1.2140127e-09, -8.977677e-10, 1.0274292e-08, 6.5348953e-09, -5.2117805e-10, -8.3820756e-10, 6.9005788e-09, 6.899254e-09, 1.3538694e-10, -7.3652023e-10, 3.4546863e-09, 6.8354673e-09, 7.216952e-10, -6.0251704e-10, 1.3999661e-10, 6.3879524e-09, 1.2110034e-09, -4.4691778e-10, -2.8669613e-09, 5.6187783e-09, 1.5846467e-09, -2.806527e-10, -5.4240217e-09, 4.602446e-09, 1.8323345e-09, -1.1421921e-10};
endpackage
`endif
