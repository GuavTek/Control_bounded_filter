`ifndef COEFFICIENTS_FX_SV_
`define COEFFICIENTS_FX_SV_
package Coefficients_Fx;
	localparam N = 4;
	localparam M = 4;
	localparam COEFF_BIAS = 48;
	localparam logic signed[63:0] Lfr[0:3] = {64'd278380577483262, 64'd278380577483262, 64'd274695218945892, 64'd274695218945892};
	localparam logic signed[63:0] Lfi[0:3] = {64'd13507030505103, - 64'd13507030505103, 64'd5413472349440, - 64'd5413472349440};
	localparam logic signed[63:0] Lbr[0:3] = {64'd278380577483262, 64'd278380577483262, 64'd274695218945892, 64'd274695218945892};
	localparam logic signed[63:0] Lbi[0:3] = {64'd13507030505103, - 64'd13507030505103, 64'd5413472349440, - 64'd5413472349440};
	localparam logic signed[63:0] Wfr[0:3] = {64'd3719944537, 64'd3719944537, - 64'd1104681121, - 64'd1104681121};
	localparam logic signed[63:0] Wfi[0:3] = {64'd152555419, - 64'd152555419, - 64'd2135740598, 64'd2135740598};
	localparam logic signed[63:0] Wbr[0:3] = {64'd3719944537, 64'd3719944537, 64'd1104681121, 64'd1104681121};
	localparam logic signed[63:0] Wbi[0:3] = {64'd152555419, - 64'd152555419, 64'd2135740598, - 64'd2135740598};
	localparam logic signed[63:0] Ffr[0:3][0:79] = '{
		'{64'd51582186096816840, 64'd5011103315704805, - 64'd561701380626195, 64'd5955993329118, 64'd53999423105038712, 64'd4657041123796227, - 64'd564755289025816, 64'd7857819238314, 64'd56238499096106752, 64'd4298618936379875, - 64'd566380727149033, 64'd9703394865811, 64'd58297472952815232, 64'd3936790712122069, - 64'd566601701445345, 64'd11489347775598, 64'd60174878023463800, 64'd3572500001736659, - 64'd565445152534737, 64'd13212516008134, 64'd61869716394208536, 64'd3206677864837182, - 64'd562940832512622, 64'd14869951625943, 64'd63381452137445600, 64'd2840240857815672, - 64'd559121177841312, 64'd16458923671137, 64'd64710003572622704, 64'd2474089096235135, - 64'd554021178222409, 64'd17976920539225, 64'd65855734577555400, 64'd2109104394973848, - 64'd547678241846547, 64'd19421651774852, 64'd66819444989881056, 64'd1746148489107903, - 64'd540132057417935, 64'd20791049296445, 64'd67602360139713424, 64'd1386061338264292, - 64'd531424453351182, 64'd22083268057958, 64'd68206119555862960, 64'd1029659516921080, - 64'd521599254536981, 64'd23296686157126, 64'd68632764889162000, 64'd677734692874472, - 64'd510702137071341, 64'd24429904400804, 64'd68884727097479536, 64'd331052195835459, - 64'd498780481340296, 64'd25481745339046, 64'd68964812937927824, - 64'd9650322138070, - 64'd485883223848305, 64'd26451251780680, 64'd68876190812551440, - 64'd343664132923856, - 64'd472060708174047, 64'd27337684804110, 64'd68622376014450832, - 64'd670310584136954, - 64'd457364535431876, 64'd28140521278033, 64'd68207215421827248, - 64'd988942155507464, - 64'd441847414611048, 64'd28859450907683, 64'd67634871687844624, - 64'd1298943419140937, - 64'd425563013157815, 64'd29494372823037, 64'd66909806974488848, - 64'd1599731903214576, - 64'd408565808157754, 64'd30045391726208},
		'{64'd51582186096781952, 64'd5011103315708102, - 64'd561701380626144, 64'd5955993329108, 64'd53999423105005552, 64'd4657041123799363, - 64'd564755289025768, 64'd7857819238304, 64'd56238499096075352, 64'd4298618936382845, - 64'd566380727148988, 64'd9703394865802, 64'd58297472952785640, 64'd3936790712124870, - 64'd566601701445303, 64'd11489347775589, 64'd60174878023436056, 64'd3572500001739287, - 64'd565445152534698, 64'd13212516008126, 64'd61869716394182680, 64'd3206677864839634, - 64'd562940832512586, 64'd14869951625935, 64'd63381452137421632, 64'd2840240857817945, - 64'd559121177841279, 64'd16458923671130, 64'd64710003572600656, 64'd2474089096237228, - 64'd554021178222378, 64'd17976920539219, 64'd65855734577535304, 64'd2109104394975759, - 64'd547678241846520, 64'd19421651774846, 64'd66819444989862912, 64'd1746148489109631, - 64'd540132057417911, 64'd20791049296440, 64'd67602360139697232, 64'd1386061338265836, - 64'd531424453351161, 64'd22083268057953, 64'd68206119555848736, 64'd1029659516922441, - 64'd521599254536963, 64'd23296686157123, 64'd68632764889149720, 64'd677734692875649, - 64'd510702137071326, 64'd24429904400801, 64'd68884727097469200, 64'd331052195836454, - 64'd498780481340284, 64'd25481745339043, 64'd68964812937919424, - 64'd9650322137257, - 64'd485883223848297, 64'd26451251780678, 64'd68876190812544960, - 64'd343664132923223, - 64'd472060708174041, 64'd27337684804109, 64'd68622376014446240, - 64'd670310584136498, - 64'd457364535431873, 64'd28140521278032, 64'd68207215421824520, - 64'd988942155507184, - 64'd441847414611048, 64'd28859450907683, 64'd67634871687843744, - 64'd1298943419140831, - 64'd425563013157818, 64'd29494372823037, 64'd66909806974489768, - 64'd1599731903214640, - 64'd408565808157760, 64'd30045391726209},
		'{- 64'd51230291296731632, - 64'd4979745320671008, 64'd540750075430615, - 64'd74242651348786, - 64'd53635973253266008, - 64'd4644905457143963, 64'd511125525001550, - 64'd71475704560060, - 64'd55877094717808200, - 64'd4321464847687858, 64'd482414340128880, - 64'd68771515801948, - 64'd57959297554849128, - 64'd4009192470127291, 64'd454600666018923, - 64'd66129690567727, - 64'd59888108183777776, - 64'd3707857601462554, 64'd427668543908287, - 64'd63549793731945, - 64'd61668937780167608, - 64'd3417230022940273, 64'd401601931135273, - 64'd61031351881953, - 64'd63307082577045232, - 64'd3137080214960943, 64'd376384720343153, - 64'd58573855575703, - 64'd64807724261133504, - 64'd2867179542118097, 64'd352000757838078, - 64'd56176761527167, - 64'd66175930459207656, - 64'd2607300428659344, 64'd328433861124088, - 64'd53839494720698, - 64'd67416655309846944, - 64'd2357216524654874, 64'd305667835637437, - 64'd51561450455693, - 64'd68534740116006152, - 64'd2116702863154401, 64'd283686490702124, - 64'd49341996322905, - 64'd69534914073970184, - 64'd1885536008608764, 64'd262473654728280, - 64'd47180474113749, - 64'd70421795074392344, - 64'd1663494196827712, 64'd242013189674693, - 64'd45076201663955, - 64'd71199890571251144, - 64'd1450357466740580, 64'd222289004796501, - 64'd43028474632921, - 64'd71873598514692880, - 64'd1245907784221772, 64'd203285069698750, - 64'd41036568220105, - 64'd72447208343856688, - 64'd1049929158238129, 64'd184985426716177, - 64'd39099738819803, - 64'd72924902035906544, - 64'd862207749570436, 64'd167374202639291, - 64'd37217225615649, - 64'd73310755207619008, - 64'd682531972356423, 64'd150435619806478, - 64'd35388252116167, - 64'd73608738265998560, - 64'd510692588697806, 64'd134154006581522, - 64'd33612027632708, - 64'd73822717604512016, - 64'd346482796569006, 64'd118513807235619, - 64'd31887748701075},
		'{- 64'd51230291296626208, - 64'd4979745320680849, 64'd540750075430448, - 64'd74242651348753, - 64'd53635973253163648, - 64'd4644905457153517, 64'd511125525001389, - 64'd71475704560028, - 64'd55877094717708872, - 64'd4321464847697130, 64'd482414340128723, - 64'd68771515801916, - 64'd57959297554752768, - 64'd4009192470136285, 64'd454600666018771, - 64'd66129690567696, - 64'd59888108183684344, - 64'd3707857601471275, 64'd427668543908139, - 64'd63549793731916, - 64'd61668937780077056, - 64'd3417230022948725, 64'd401601931135130, - 64'd61031351881925, - 64'd63307082576957520, - 64'd3137080214969132, 64'd376384720343014, - 64'd58573855575676, - 64'd64807724261048560, - 64'd2867179542126026, 64'd352000757837944, - 64'd56176761527141, - 64'd66175930459125448, - 64'd2607300428667019, 64'd328433861123959, - 64'd53839494720672, - 64'd67416655309767400, - 64'd2357216524662300, 64'd305667835637311, - 64'd51561450455668, - 64'd68534740115929232, - 64'd2116702863161581, 64'd283686490702003, - 64'd49341996322881, - 64'd69534914073895848, - 64'd1885536008615703, 64'd262473654728163, - 64'd47180474113726, - 64'd70421795074320528, - 64'd1663494196834416, 64'd242013189674580, - 64'd45076201663933, - 64'd71199890571181800, - 64'd1450357466747053, 64'd222289004796392, - 64'd43028474632899, - 64'd71873598514625968, - 64'd1245907784228020, 64'd203285069698645, - 64'd41036568220084, - 64'd72447208343792128, - 64'd1049929158244155, 64'd184985426716076, - 64'd39099738819783, - 64'd72924902035844320, - 64'd862207749576246, 64'd167374202639194, - 64'd37217225615629, - 64'd73310755207559056, - 64'd682531972362020, 64'd150435619806384, - 64'd35388252116148, - 64'd73608738265940832, - 64'd510692588703196, 64'd134154006581431, - 64'd33612027632690, - 64'd73822717604456448, - 64'd346482796574194, 64'd118513807235532, - 64'd31887748701058}};
	localparam logic signed[63:0] Ffi[0:3][0:79] = '{
		'{- 64'd62190398332284048, 64'd6230332637606097, 64'd192324072483146, - 64'd40996918193475, - 64'd59031452936600264, 64'd6402305256326630, 64'd163255608778863, - 64'd40260410039214, - 64'd55791240438299936, 64'd6555397046536509, 64'd134360162933161, - 64'd39440736515934, - 64'd52479203592061040, 64'd6689606353484126, 64'd105704380320668, - 64'd38541511163769, - 64'd49104774491139680, 64'd6804977317853832, 64'd77353021660942, - 64'd37566469629123, - 64'd45677351916584496, 64'd6901598872870764, 64'd49368842936556, - 64'd36519458222243, - 64'd42206279210313192, 64'd6979603652467820, 64'd21812482519020, - 64'd35404422430442, - 64'd38700822715428976, 64'd7039166814900830, - 64'd5257644364900, - 64'd34225395415677, - 64'd35170150824931108, 64'd7080504786317119, - 64'd31785443714318, - 64'd32986486524670, - 64'd31623313677694240, 64'd7103873928888477, - 64'd57717233290888, - 64'd31691869839176, - 64'd28069223538262032, 64'd7109569138212226, - 64'd83001825539176, - 64'd30345772793346, - 64'd24516635894628184, 64'd7097922374763421, - 64'd107590602838786, - 64'd28952464884485, - 64'd20974131305769588, 64'd7069301134247510, - 64'd131437585055862, - 64'd27516246502709, - 64'd17450098028257504, 64'd7024106861755984, - 64'd154499489380911, - 64'd26041437904274, - 64'd13952715448811096, 64'd6962773314667836, - 64'd176735782458836, - 64'd24532368352469, - 64'd10489938347178780, 64'd6885764879267162, - 64'd198108724835619, - 64'd22993365449127, - 64'd7069482011243008, 64'd6793574846062164, - 64'd218583407764256, - 64'd21428744678871, - 64'd3698808223751144, 64'd6686723648793412, - 64'd238127782430210, - 64'd19842799187279, - 64'd385112137582196, 64'd6565757072109603, - 64'd256712681673870, - 64'd18239789813167, 64'd2864689946024472, 64'd6431244432867604, - 64'd274311834304139, - 64'd16623935394169},
		'{64'd62190398332311936, - 64'd6230332637608698, - 64'd192324072483193, 64'd40996918193485, 64'd59031452936629520, - 64'd6402305256329361, - 64'd163255608778913, 64'd40260410039224, 64'd55791240438330464, - 64'd6555397046539360, - 64'd134360162933213, 64'd39440736515945, 64'd52479203592092736, - 64'd6689606353487088, - 64'd105704380320721, 64'd38541511163780, 64'd49104774491172456, - 64'd6804977317856896, - 64'd77353021660996, 64'd37566469629134, 64'd45677351916618240, - 64'd6901598872873920, - 64'd49368842936611, 64'd36519458222254, 64'd42206279210347800, - 64'd6979603652471059, - 64'd21812482519077, 64'd35404422430454, 64'd38700822715464344, - 64'd7039166814904143, 64'd5257644364842, 64'd34225395415688, 64'd35170150824967148, - 64'd7080504786320496, 64'd31785443714260, 64'd32986486524682, 64'd31623313677730856, - 64'd7103873928891909, 64'd57717233290828, 64'd31691869839188, 64'd28069223538299116, - 64'd7109569138215704, 64'd83001825539116, 64'd30345772793358, 64'd24516635894665640, - 64'd7097922374766934, 64'd107590602838726, 64'd28952464884497, 64'd20974131305807312, - 64'd7069301134251049, 64'd131437585055802, 64'd27516246502721, 64'd17450098028295404, - 64'd7024106861759542, 64'd154499489380850, 64'd26041437904286, 64'd13952715448849076, - 64'd6962773314671402, 64'd176735782458775, 64'd24532368352481, 64'd10489938347216740, - 64'd6885764879270728, 64'd198108724835559, 64'd22993365449139, 64'd7069482011280864, - 64'd6793574846065721, 64'd218583407764196, 64'd21428744678883, 64'd3698808223788804, - 64'd6686723648796952, 64'd238127782430150, 64'd19842799187291, 64'd385112137619572, - 64'd6565757072113116, 64'd256712681673812, 64'd18239789813179, - 64'd2864689945987468, - 64'd6431244432871084, 64'd274311834304082, 64'd16623935394181},
		'{64'd189244198874480864, - 64'd11173526320859200, 64'd863108706904317, - 64'd50887687823156, 64'd183700673796767296, - 64'd11000167790722104, 64'd852719391270143, - 64'd51089852662961, 64'd178244405727557888, - 64'd10824545053978236, 64'd842010563605728, - 64'd51233932699752, 64'd172876457860091936, - 64'd10646931883877146, 64'd831007486168611, - 64'd51322533990261, 64'd167597759271707968, - 64'd10467591016280584, 64'd819734507808407, - 64'd51358192232975, 64'd162409110374531552, - 64'd10286774421268872, 64'd808215083968045, - 64'd51343373681628, 64'd157311188231003232, - 64'd10104723572149220, 64'd796471796589263, - 64'd51280476081521, 64'd152304551735580256, - 64'd9921669711733166, 64'd784526373907983, - 64'd51171829626718, 64'd147389646664007872, - 64'd9737834115759036, 64'd772399710125948, - 64'd51019697936218, 64'd142566810591617232, - 64'd9553428353344048, 64'd760111884945779, - 64'd50826279047275, 64'd137836277682162752, - 64'd9368654544358890, 64'd747682182957348, - 64'd50593706424120, 64'd133198183348761952, - 64'd9183705613625504, 64'd735129112864062, - 64'd50324049980397, 64'd128652568788549888, - 64'd8998765541846701, 64'd722470426538354, - 64'd50019317113685, 64'd124199385392703584, - 64'd8814009613183452, 64'd709723137896350, - 64'd49681453750570, 64'd119838499033531904, - 64'd8629604659403012, 64'd696903541582309, - 64'd49312345400761, 64'd115569694230363168, - 64'd8445709300527816, 64'd684027231454067, - 64'd48913818218825, 64'd111392678195997040, - 64'd8262474181921818, 64'd671109118861341, - 64'd48487640072178, 64'd107307084765515040, - 64'd8080042207757172, 64'd658163450709275, - 64'd48035521614017, 64'd103312478209274096, - 64'd7898548770810504, 64'd645203827300241, - 64'd47559117359940, 64'd99408356931928416, - 64'd7718121978543659, 64'd632243219947395, - 64'd47060026767058},
		'{- 64'd189244198874508576, 64'd11173526320861784, - 64'd863108706904270, 64'd50887687823147, - 64'd183700673796796384, 64'd11000167790724812, - 64'd852719391270094, 64'd51089852662951, - 64'd178244405727588192, 64'd10824545053981066, - 64'd842010563605678, 64'd51233932699742, - 64'd172876457860123456, 64'd10646931883880084, - 64'd831007486168558, 64'd51322533990250, - 64'd167597759271740608, 64'd10467591016283628, - 64'd819734507808353, 64'd51358192232964, - 64'd162409110374565152, 64'd10286774421272006, - 64'd808215083967989, 64'd51343373681617, - 64'd157311188231037792, 64'd10104723572152444, - 64'd796471796589206, 64'd51280476081509, - 64'd152304551735615648, 64'd9921669711736470, - 64'd784526373907925, 64'd51171829626706, - 64'd147389646664044096, 64'd9737834115762410, - 64'd772399710125888, 64'd51019697936206, - 64'd142566810591654144, 64'd9553428353347490, - 64'd760111884945718, 64'd50826279047263, - 64'd137836277682200304, 64'd9368654544362392, - 64'd747682182957286, 64'd50593706424108, - 64'd133198183348800064, 64'd9183705613629060, - 64'd735129112863999, 64'd50324049980384, - 64'd128652568788588528, 64'd8998765541850306, - 64'd722470426538291, 64'd50019317113672, - 64'd124199385392742656, 64'd8814009613187097, - 64'd709723137896286, 64'd49681453750558, - 64'd119838499033571376, 64'd8629604659406695, - 64'd696903541582244, 64'd49312345400748, - 64'd115569694230402960, 64'd8445709300531530, - 64'd684027231454002, 64'd48913818218812, - 64'd111392678196037120, 64'd8262474181925558, - 64'd671109118861276, 64'd48487640072165, - 64'd107307084765555360, 64'd8080042207760935, - 64'd658163450709210, 64'd48035521614004, - 64'd103312478209314576, 64'd7898548770814283, - 64'd645203827300175, 64'd47559117359927, - 64'd99408356931969056, 64'd7718121978547451, - 64'd632243219947328, 64'd47060026767044}};
	localparam logic signed[63:0] Fbr[0:3][0:79] = '{
		'{64'd51582186096816840, - 64'd5011103315704805, - 64'd561701380626195, - 64'd5955993329118, 64'd53999423105038712, - 64'd4657041123796227, - 64'd564755289025816, - 64'd7857819238314, 64'd56238499096106752, - 64'd4298618936379875, - 64'd566380727149033, - 64'd9703394865811, 64'd58297472952815232, - 64'd3936790712122069, - 64'd566601701445345, - 64'd11489347775598, 64'd60174878023463800, - 64'd3572500001736659, - 64'd565445152534737, - 64'd13212516008134, 64'd61869716394208536, - 64'd3206677864837182, - 64'd562940832512622, - 64'd14869951625943, 64'd63381452137445600, - 64'd2840240857815672, - 64'd559121177841312, - 64'd16458923671137, 64'd64710003572622704, - 64'd2474089096235135, - 64'd554021178222409, - 64'd17976920539225, 64'd65855734577555400, - 64'd2109104394973848, - 64'd547678241846547, - 64'd19421651774852, 64'd66819444989881056, - 64'd1746148489107903, - 64'd540132057417935, - 64'd20791049296445, 64'd67602360139713424, - 64'd1386061338264292, - 64'd531424453351182, - 64'd22083268057958, 64'd68206119555862960, - 64'd1029659516921080, - 64'd521599254536981, - 64'd23296686157126, 64'd68632764889162000, - 64'd677734692874472, - 64'd510702137071341, - 64'd24429904400804, 64'd68884727097479536, - 64'd331052195835459, - 64'd498780481340296, - 64'd25481745339046, 64'd68964812937927824, 64'd9650322138070, - 64'd485883223848305, - 64'd26451251780680, 64'd68876190812551440, 64'd343664132923856, - 64'd472060708174047, - 64'd27337684804110, 64'd68622376014450832, 64'd670310584136954, - 64'd457364535431876, - 64'd28140521278033, 64'd68207215421827248, 64'd988942155507464, - 64'd441847414611048, - 64'd28859450907683, 64'd67634871687844624, 64'd1298943419140937, - 64'd425563013157815, - 64'd29494372823037, 64'd66909806974488848, 64'd1599731903214576, - 64'd408565808157754, - 64'd30045391726208},
		'{64'd51582186096781952, - 64'd5011103315708102, - 64'd561701380626144, - 64'd5955993329108, 64'd53999423105005552, - 64'd4657041123799363, - 64'd564755289025768, - 64'd7857819238304, 64'd56238499096075352, - 64'd4298618936382845, - 64'd566380727148988, - 64'd9703394865802, 64'd58297472952785640, - 64'd3936790712124870, - 64'd566601701445303, - 64'd11489347775589, 64'd60174878023436056, - 64'd3572500001739287, - 64'd565445152534698, - 64'd13212516008126, 64'd61869716394182680, - 64'd3206677864839634, - 64'd562940832512586, - 64'd14869951625935, 64'd63381452137421632, - 64'd2840240857817945, - 64'd559121177841279, - 64'd16458923671130, 64'd64710003572600656, - 64'd2474089096237228, - 64'd554021178222378, - 64'd17976920539219, 64'd65855734577535304, - 64'd2109104394975759, - 64'd547678241846520, - 64'd19421651774846, 64'd66819444989862912, - 64'd1746148489109631, - 64'd540132057417911, - 64'd20791049296440, 64'd67602360139697232, - 64'd1386061338265836, - 64'd531424453351161, - 64'd22083268057953, 64'd68206119555848736, - 64'd1029659516922441, - 64'd521599254536963, - 64'd23296686157123, 64'd68632764889149720, - 64'd677734692875649, - 64'd510702137071326, - 64'd24429904400801, 64'd68884727097469200, - 64'd331052195836454, - 64'd498780481340284, - 64'd25481745339043, 64'd68964812937919424, 64'd9650322137257, - 64'd485883223848297, - 64'd26451251780678, 64'd68876190812544960, 64'd343664132923223, - 64'd472060708174041, - 64'd27337684804109, 64'd68622376014446240, 64'd670310584136498, - 64'd457364535431873, - 64'd28140521278032, 64'd68207215421824520, 64'd988942155507184, - 64'd441847414611048, - 64'd28859450907683, 64'd67634871687843744, 64'd1298943419140831, - 64'd425563013157818, - 64'd29494372823037, 64'd66909806974489768, 64'd1599731903214640, - 64'd408565808157760, - 64'd30045391726209},
		'{64'd51230291296731632, - 64'd4979745320671008, - 64'd540750075430615, - 64'd74242651348786, 64'd53635973253266008, - 64'd4644905457143963, - 64'd511125525001550, - 64'd71475704560060, 64'd55877094717808200, - 64'd4321464847687858, - 64'd482414340128880, - 64'd68771515801948, 64'd57959297554849128, - 64'd4009192470127291, - 64'd454600666018923, - 64'd66129690567727, 64'd59888108183777776, - 64'd3707857601462554, - 64'd427668543908287, - 64'd63549793731945, 64'd61668937780167608, - 64'd3417230022940273, - 64'd401601931135273, - 64'd61031351881953, 64'd63307082577045232, - 64'd3137080214960943, - 64'd376384720343153, - 64'd58573855575703, 64'd64807724261133504, - 64'd2867179542118097, - 64'd352000757838078, - 64'd56176761527167, 64'd66175930459207656, - 64'd2607300428659344, - 64'd328433861124088, - 64'd53839494720698, 64'd67416655309846944, - 64'd2357216524654874, - 64'd305667835637437, - 64'd51561450455693, 64'd68534740116006152, - 64'd2116702863154401, - 64'd283686490702124, - 64'd49341996322905, 64'd69534914073970184, - 64'd1885536008608764, - 64'd262473654728280, - 64'd47180474113749, 64'd70421795074392344, - 64'd1663494196827712, - 64'd242013189674693, - 64'd45076201663955, 64'd71199890571251144, - 64'd1450357466740580, - 64'd222289004796501, - 64'd43028474632921, 64'd71873598514692880, - 64'd1245907784221772, - 64'd203285069698750, - 64'd41036568220105, 64'd72447208343856688, - 64'd1049929158238129, - 64'd184985426716177, - 64'd39099738819803, 64'd72924902035906544, - 64'd862207749570436, - 64'd167374202639291, - 64'd37217225615649, 64'd73310755207619008, - 64'd682531972356423, - 64'd150435619806478, - 64'd35388252116167, 64'd73608738265998560, - 64'd510692588697806, - 64'd134154006581522, - 64'd33612027632708, 64'd73822717604512016, - 64'd346482796569006, - 64'd118513807235619, - 64'd31887748701075},
		'{64'd51230291296626208, - 64'd4979745320680849, - 64'd540750075430448, - 64'd74242651348753, 64'd53635973253163648, - 64'd4644905457153517, - 64'd511125525001389, - 64'd71475704560028, 64'd55877094717708872, - 64'd4321464847697130, - 64'd482414340128723, - 64'd68771515801916, 64'd57959297554752768, - 64'd4009192470136285, - 64'd454600666018771, - 64'd66129690567696, 64'd59888108183684344, - 64'd3707857601471275, - 64'd427668543908139, - 64'd63549793731916, 64'd61668937780077056, - 64'd3417230022948725, - 64'd401601931135130, - 64'd61031351881925, 64'd63307082576957520, - 64'd3137080214969132, - 64'd376384720343014, - 64'd58573855575676, 64'd64807724261048560, - 64'd2867179542126026, - 64'd352000757837944, - 64'd56176761527141, 64'd66175930459125448, - 64'd2607300428667019, - 64'd328433861123959, - 64'd53839494720672, 64'd67416655309767400, - 64'd2357216524662300, - 64'd305667835637311, - 64'd51561450455668, 64'd68534740115929232, - 64'd2116702863161581, - 64'd283686490702003, - 64'd49341996322881, 64'd69534914073895848, - 64'd1885536008615703, - 64'd262473654728163, - 64'd47180474113726, 64'd70421795074320528, - 64'd1663494196834416, - 64'd242013189674580, - 64'd45076201663933, 64'd71199890571181800, - 64'd1450357466747053, - 64'd222289004796392, - 64'd43028474632899, 64'd71873598514625968, - 64'd1245907784228020, - 64'd203285069698645, - 64'd41036568220084, 64'd72447208343792128, - 64'd1049929158244155, - 64'd184985426716076, - 64'd39099738819783, 64'd72924902035844320, - 64'd862207749576246, - 64'd167374202639194, - 64'd37217225615629, 64'd73310755207559056, - 64'd682531972362020, - 64'd150435619806384, - 64'd35388252116148, 64'd73608738265940832, - 64'd510692588703196, - 64'd134154006581431, - 64'd33612027632690, 64'd73822717604456448, - 64'd346482796574194, - 64'd118513807235532, - 64'd31887748701058}};
	localparam logic signed[63:0] Fbi[0:3][0:79] = '{
		'{- 64'd62190398332284048, - 64'd6230332637606097, 64'd192324072483146, 64'd40996918193475, - 64'd59031452936600264, - 64'd6402305256326630, 64'd163255608778863, 64'd40260410039214, - 64'd55791240438299936, - 64'd6555397046536509, 64'd134360162933161, 64'd39440736515934, - 64'd52479203592061040, - 64'd6689606353484126, 64'd105704380320668, 64'd38541511163769, - 64'd49104774491139680, - 64'd6804977317853832, 64'd77353021660942, 64'd37566469629123, - 64'd45677351916584496, - 64'd6901598872870764, 64'd49368842936556, 64'd36519458222243, - 64'd42206279210313192, - 64'd6979603652467820, 64'd21812482519020, 64'd35404422430442, - 64'd38700822715428976, - 64'd7039166814900830, - 64'd5257644364900, 64'd34225395415677, - 64'd35170150824931108, - 64'd7080504786317119, - 64'd31785443714318, 64'd32986486524670, - 64'd31623313677694240, - 64'd7103873928888477, - 64'd57717233290888, 64'd31691869839176, - 64'd28069223538262032, - 64'd7109569138212226, - 64'd83001825539176, 64'd30345772793346, - 64'd24516635894628184, - 64'd7097922374763421, - 64'd107590602838786, 64'd28952464884485, - 64'd20974131305769588, - 64'd7069301134247510, - 64'd131437585055862, 64'd27516246502709, - 64'd17450098028257504, - 64'd7024106861755984, - 64'd154499489380911, 64'd26041437904274, - 64'd13952715448811096, - 64'd6962773314667836, - 64'd176735782458836, 64'd24532368352469, - 64'd10489938347178780, - 64'd6885764879267162, - 64'd198108724835619, 64'd22993365449127, - 64'd7069482011243008, - 64'd6793574846062164, - 64'd218583407764256, 64'd21428744678871, - 64'd3698808223751144, - 64'd6686723648793412, - 64'd238127782430210, 64'd19842799187279, - 64'd385112137582196, - 64'd6565757072109603, - 64'd256712681673870, 64'd18239789813167, 64'd2864689946024472, - 64'd6431244432867604, - 64'd274311834304139, 64'd16623935394169},
		'{64'd62190398332311936, 64'd6230332637608698, - 64'd192324072483193, - 64'd40996918193485, 64'd59031452936629520, 64'd6402305256329361, - 64'd163255608778913, - 64'd40260410039224, 64'd55791240438330464, 64'd6555397046539360, - 64'd134360162933213, - 64'd39440736515945, 64'd52479203592092736, 64'd6689606353487088, - 64'd105704380320721, - 64'd38541511163780, 64'd49104774491172456, 64'd6804977317856896, - 64'd77353021660996, - 64'd37566469629134, 64'd45677351916618240, 64'd6901598872873920, - 64'd49368842936611, - 64'd36519458222254, 64'd42206279210347800, 64'd6979603652471059, - 64'd21812482519077, - 64'd35404422430454, 64'd38700822715464344, 64'd7039166814904143, 64'd5257644364842, - 64'd34225395415688, 64'd35170150824967148, 64'd7080504786320496, 64'd31785443714260, - 64'd32986486524682, 64'd31623313677730856, 64'd7103873928891909, 64'd57717233290828, - 64'd31691869839188, 64'd28069223538299116, 64'd7109569138215704, 64'd83001825539116, - 64'd30345772793358, 64'd24516635894665640, 64'd7097922374766934, 64'd107590602838726, - 64'd28952464884497, 64'd20974131305807312, 64'd7069301134251049, 64'd131437585055802, - 64'd27516246502721, 64'd17450098028295404, 64'd7024106861759542, 64'd154499489380850, - 64'd26041437904286, 64'd13952715448849076, 64'd6962773314671402, 64'd176735782458775, - 64'd24532368352481, 64'd10489938347216740, 64'd6885764879270728, 64'd198108724835559, - 64'd22993365449139, 64'd7069482011280864, 64'd6793574846065721, 64'd218583407764196, - 64'd21428744678883, 64'd3698808223788804, 64'd6686723648796952, 64'd238127782430150, - 64'd19842799187291, 64'd385112137619572, 64'd6565757072113116, 64'd256712681673812, - 64'd18239789813179, - 64'd2864689945987468, 64'd6431244432871084, 64'd274311834304082, - 64'd16623935394181},
		'{- 64'd189244198874480864, - 64'd11173526320859200, - 64'd863108706904317, - 64'd50887687823156, - 64'd183700673796767296, - 64'd11000167790722104, - 64'd852719391270143, - 64'd51089852662961, - 64'd178244405727557888, - 64'd10824545053978236, - 64'd842010563605728, - 64'd51233932699752, - 64'd172876457860091936, - 64'd10646931883877146, - 64'd831007486168611, - 64'd51322533990261, - 64'd167597759271707968, - 64'd10467591016280584, - 64'd819734507808407, - 64'd51358192232975, - 64'd162409110374531552, - 64'd10286774421268872, - 64'd808215083968045, - 64'd51343373681628, - 64'd157311188231003232, - 64'd10104723572149220, - 64'd796471796589263, - 64'd51280476081521, - 64'd152304551735580256, - 64'd9921669711733166, - 64'd784526373907983, - 64'd51171829626718, - 64'd147389646664007872, - 64'd9737834115759036, - 64'd772399710125948, - 64'd51019697936218, - 64'd142566810591617232, - 64'd9553428353344048, - 64'd760111884945779, - 64'd50826279047275, - 64'd137836277682162752, - 64'd9368654544358890, - 64'd747682182957348, - 64'd50593706424120, - 64'd133198183348761952, - 64'd9183705613625504, - 64'd735129112864062, - 64'd50324049980397, - 64'd128652568788549888, - 64'd8998765541846701, - 64'd722470426538354, - 64'd50019317113685, - 64'd124199385392703584, - 64'd8814009613183452, - 64'd709723137896350, - 64'd49681453750570, - 64'd119838499033531904, - 64'd8629604659403012, - 64'd696903541582309, - 64'd49312345400761, - 64'd115569694230363168, - 64'd8445709300527816, - 64'd684027231454067, - 64'd48913818218825, - 64'd111392678195997040, - 64'd8262474181921818, - 64'd671109118861341, - 64'd48487640072178, - 64'd107307084765515040, - 64'd8080042207757172, - 64'd658163450709275, - 64'd48035521614017, - 64'd103312478209274096, - 64'd7898548770810504, - 64'd645203827300241, - 64'd47559117359940, - 64'd99408356931928416, - 64'd7718121978543659, - 64'd632243219947395, - 64'd47060026767058},
		'{64'd189244198874508576, 64'd11173526320861784, 64'd863108706904270, 64'd50887687823147, 64'd183700673796796384, 64'd11000167790724812, 64'd852719391270094, 64'd51089852662951, 64'd178244405727588192, 64'd10824545053981066, 64'd842010563605678, 64'd51233932699742, 64'd172876457860123456, 64'd10646931883880084, 64'd831007486168558, 64'd51322533990250, 64'd167597759271740608, 64'd10467591016283628, 64'd819734507808353, 64'd51358192232964, 64'd162409110374565152, 64'd10286774421272006, 64'd808215083967989, 64'd51343373681617, 64'd157311188231037792, 64'd10104723572152444, 64'd796471796589206, 64'd51280476081509, 64'd152304551735615648, 64'd9921669711736470, 64'd784526373907925, 64'd51171829626706, 64'd147389646664044096, 64'd9737834115762410, 64'd772399710125888, 64'd51019697936206, 64'd142566810591654144, 64'd9553428353347490, 64'd760111884945718, 64'd50826279047263, 64'd137836277682200304, 64'd9368654544362392, 64'd747682182957286, 64'd50593706424108, 64'd133198183348800064, 64'd9183705613629060, 64'd735129112863999, 64'd50324049980384, 64'd128652568788588528, 64'd8998765541850306, 64'd722470426538291, 64'd50019317113672, 64'd124199385392742656, 64'd8814009613187097, 64'd709723137896286, 64'd49681453750558, 64'd119838499033571376, 64'd8629604659406695, 64'd696903541582244, 64'd49312345400748, 64'd115569694230402960, 64'd8445709300531530, 64'd684027231454002, 64'd48913818218812, 64'd111392678196037120, 64'd8262474181925558, 64'd671109118861276, 64'd48487640072165, 64'd107307084765555360, 64'd8080042207760935, 64'd658163450709210, 64'd48035521614004, 64'd103312478209314576, 64'd7898548770814283, 64'd645203827300175, 64'd47559117359927, 64'd99408356931969056, 64'd7718121978547451, 64'd632243219947328, 64'd47060026767044}};
	localparam logic signed[63:0] hf[0:1199] = {64'd4704787496960, - 64'd4776038912, - 64'd6201745920, 64'd12376386, 64'd4700013330432, - 64'd14318410752, - 64'd6176088576, 64'd37060376, 64'd4690473910272, - 64'd23831724032, - 64'd6124879360, 64'd61541484, 64'd4676189683712, - 64'd33296730112, - 64'd6048317440, 64'd85691840, 64'd4657188438016, - 64'd42694332416, - 64'd5946690560, 64'd109390016, 64'd4633509494784, - 64'd52005650432, - 64'd5820371456, 64'd132521128, 64'd4605200039936, - 64'd61212069888, - 64'd5669813760, 64'd154976880, 64'd4572317745152, - 64'd70295289856, - 64'd5495548928, 64'd176655632, 64'd4534928146432, - 64'd79237382144, - 64'd5298182656, 64'd197462448, 64'd4493106741248, - 64'd88020836352, - 64'd5078390272, 64'd217309056, 64'd4446936891392, - 64'd96628596736, - 64'd4836913152, 64'd236113952, 64'd4396510085120, - 64'd105044131840, - 64'd4574555136, 64'd253802304, 64'd4341927247872, - 64'd113251434496, - 64'd4292176128, 64'd270305984, 64'd4283295858688, - 64'd121235111936, - 64'd3990691840, 64'd285563488, 64'd4220731785216, - 64'd128980369408, - 64'd3671066112, 64'd299519904, 64'd4154357710848, - 64'd136473083904, - 64'd3334309120, 64'd312126848, 64'd4084303134720, - 64'd143699820544, - 64'd2981470976, 64'd323342368, 64'd4010704109568, - 64'd150647848960, - 64'd2613640448, 64'd333130880, 64'd3933703503872, - 64'd157305192448, - 64'd2231937536, 64'd341463008, 64'd3853449166848, - 64'd163660644352, - 64'd1837512192, 64'd348315488, 64'd3770094977024, - 64'd169703784448, - 64'd1431538176, 64'd353671104, 64'd3683799007232, - 64'd175424978944, - 64'd1015210240, 64'd357518464, 64'd3594725097472, - 64'd180815462400, - 64'd589739520, 64'd359851872, 64'd3503039971328, - 64'd185867239424, - 64'd156349744, 64'd360671232, 64'd3408915333120, - 64'd190573232128, 64'd283726752, 64'd359981728, 64'd3312525508608, - 64'd194927149056, 64'd729252672, 64'd357793824, 64'd3214047707136, - 64'd198923616256, 64'd1178989696, 64'd354122944, 64'd3113662283776, - 64'd202558095360, 64'd1631701888, 64'd348989408, 64'd3011550642176, - 64'd205826899968, 64'd2086159488, 64'd342418112, 64'd2907896545280, - 64'd208727244800, 64'd2541142016, 64'd334438336, 64'd2802885066752, - 64'd211257163776, 64'd2995442432, 64'd325083616, 64'd2696701280256, - 64'd213415575552, 64'd3447869184, 64'd314391488, 64'd2589531570176, - 64'd215202234368, 64'd3897250048, 64'd302403232, 64'd2481561010176, - 64'd216617730048, 64'd4342434816, 64'd289163680, 64'd2372975460352, - 64'd217663455232, 64'd4782299136, 64'd274721024, 64'd2263958683648, - 64'd218341638144, 64'd5215745024, 64'd259126464, 64'd2154694443008, - 64'd218655309824, 64'd5641705984, 64'd242434144, 64'd2045363617792, - 64'd218608222208, 64'd6059147776, 64'd224700832, 64'd1936145645568, - 64'd218204946432, 64'd6467070976, 64'd205985664, 64'd1827217211392, - 64'd217450758144, 64'd6864514560, 64'd186349936, 64'd1718752378880, - 64'd216351637504, 64'd7250554880, 64'd165856928, 64'd1610921934848, - 64'd214914269184, 64'd7624310784, 64'd144571552, 64'd1503893258240, - 64'd213145993216, 64'd7984943616, 64'd122560264, 64'd1397829795840, - 64'd211054772224, 64'd8331659264, 64'd99890704, 64'd1292890800128, - 64'd208649191424, 64'd8663708672, 64'd76631560, 64'd1189231460352, - 64'd205938409472, 64'd8980389888, 64'd52852316, 64'd1087001722880, - 64'd202932142080, 64'd9281050624, 64'd28623022, 64'd986346881024, - 64'd199640612864, 64'd9565084672, 64'd4014100, 64'd887406854144, - 64'd196074520576, 64'd9831939072, - 64'd20903884, 64'd790316253184, - 64'd192245039104, 64'd10081110016, - 64'd46060420, 64'd695203790848, - 64'd188163735552, 64'd10312142848, - 64'd71385240, 64'd602192478208, - 64'd183842586624, 64'd10524638208, - 64'd96808552, 64'd511399165952, - 64'd179293913088, 64'd10718244864, - 64'd122261184, 64'd422934413312, - 64'd174530363392, 64'd10892664832, - 64'd147674800, 64'd336902488064, - 64'd169564848128, 64'd11047652352, - 64'd172982048, 64'd253401055232, - 64'd164410523648, 64'd11183011840, - 64'd198116768, 64'd172521209856, - 64'd159080792064, 64'd11298598912, - 64'd223014128, 64'd94347255808, - 64'd153589219328, 64'd11394321408, - 64'd247610784, 64'd18956701696, - 64'd147949502464, 64'd11470135296, - 64'd271845024, - 64'd53579837440, - 64'd142175469568, 64'd11526046720, - 64'd295656928, - 64'd123198676992, - 64'd136281006080, 64'd11562112000, - 64'd318988480, - 64'd189843079168, - 64'd130280062976, 64'd11578433536, - 64'd341783712, - 64'd253463298048, - 64'd124186583040, 64'd11575159808, - 64'd363988800, - 64'd314016530432, - 64'd118014500864, 64'd11552485376, - 64'd385552160, - 64'd371466993664, - 64'd111777677312, 64'd11510649856, - 64'd406424608, - 64'd425785720832, - 64'd105489899520, 64'd11449936896, - 64'd426559392, - 64'd476950659072, - 64'd99164839936, 64'd11370668032, - 64'd445912288, - 64'd524946571264, - 64'd92816015360, 64'd11273207808, - 64'd464441728, - 64'd569764937728, - 64'd86456786944, 64'd11157959680, - 64'd482108768, - 64'd611403759616, - 64'd80100278272, 64'd11025362944, - 64'd498877216, - 64'd649867821056, - 64'd73759424512, 64'd10875890688, - 64'd514713696, - 64'd685167935488, - 64'd67446861824, 64'd10710052864, - 64'd529587616, - 64'd717321404416, - 64'd61174980608, 64'd10528389120, - 64'd543471232, - 64'd746351689728, - 64'd54955843584, 64'd10331468800, - 64'd556339776, - 64'd772288020480, - 64'd48801189888, 64'd10119888896, - 64'd568171200, - 64'd795165523968, - 64'd42722418688, 64'd9894274048, - 64'd578946624, - 64'd815024898048, - 64'd36730548224, 64'd9655272448, - 64'd588649792, - 64'd831912280064, - 64'd30836209664, 64'd9403553792, - 64'd597267584, - 64'd845879050240, - 64'd25049632768, 64'd9139807232, - 64'd604789568, - 64'd856981504000, - 64'd19380617216, 64'd8864742400, - 64'd611208448, - 64'd865280786432, - 64'd13838529536, 64'd8579081728, - 64'd616519488, - 64'd870842630144, - 64'd8432279040, 64'd8283564544, - 64'd620720832, - 64'd873737093120, - 64'd3170313216, 64'd7978940416, - 64'd623813568, - 64'd874038362112, 64'd1939399552, 64'd7665970176, - 64'd625801280, - 64'd871824359424, 64'd6889375744, 64'd7345421312, - 64'd626690240, - 64'd867176742912, 64'd11672628224, 64'd7018067968, - 64'd626489408, - 64'd860180578304, 64'd16282670080, 64'd6684688384, - 64'd625210304, - 64'd850923945984, 64'd20713525248, 64'd6346062848, - 64'd622866752, - 64'd839497809920, 64'd24959727616, 64'd6002970624, - 64'd619475072, - 64'd825995821056, 64'd29016330240, 64'd5656191488, - 64'd615053952, - 64'd810513793024, 64'd32878905344, 64'd5306499072, - 64'd609624128, - 64'd793149898752, 64'd36543541248, 64'd4954663936, - 64'd603208640, - 64'd774003818496, 64'd40006840320, 64'd4601447424, - 64'd595832512, - 64'd753177067520, 64'd43265937408, 64'd4247603456, - 64'd587522624, - 64'd730772340736, 64'd46318465024, 64'd3893874944, - 64'd578307904, - 64'd706893316096, 64'd49162575872, 64'd3540992256, - 64'd568218752, - 64'd681644720128, 64'd51796918272, 64'd3189672704, - 64'd557287488, - 64'd655131541504, 64'd54220648448, 64'd2840618240, - 64'd545547776, - 64'd627459227648, 64'd56433414144, 64'd2494514432, - 64'd533034752, - 64'd598733291520, 64'd58435334144, 64'd2152028160, - 64'd519784928, - 64'd569058918400, 64'd60227010560, 64'd1813808128, - 64'd505835904, - 64'd538541129728, 64'd61809512448, 64'd1480481920, - 64'd491226464, - 64'd507284029440, 64'd63184347136, 64'd1152655872, - 64'd475996352, - 64'd475391066112, 64'd64353472512, 64'd830913536, - 64'd460186112, - 64'd442964475904, 64'd65319268352, 64'd515814912, - 64'd443837152, - 64'd410105217024, 64'd66084532224, 64'd207895440, - 64'd426991392, - 64'd376912838656, 64'd66652459008, - 64'd92334792, - 64'd409691392, - 64'd343485054976, 64'd67026620416, - 64'd384391904, - 64'd391980032, - 64'd309917843456, 64'd67210969088, - 64'd667818816, - 64'd373900512, - 64'd276305018880, 64'd67209797632, - 64'd942185920, - 64'd355496224, - 64'd242738216960, 64'd67027738624, - 64'd1207091584, - 64'd336810688, - 64'd209306615808, 64'd66669740032, - 64'd1462162688, - 64'd317887360, - 64'd176096935936, 64'd66141057024, - 64'd1707054720, - 64'd298769568, - 64'd143193096192, 64'd65447219200, - 64'd1941452544, - 64'd279500384, - 64'd110676279296, 64'd64594018304, - 64'd2165070336, - 64'd260122560, - 64'd78624645120, 64'd63587500032, - 64'd2377651712, - 64'd240678480, - 64'd47113297920, 64'd62433927168, - 64'd2578969600, - 64'd221209920, - 64'd16214159360, 64'd61139771392, - 64'd2768827136, - 64'd201758064, 64'd14004141056, 64'd59711692800, - 64'd2947056640, - 64'd182363424, 64'd43476340736, 64'd58156523520, - 64'd3113519360, - 64'd163065696, 64'd72140636160, 64'd56481234944, - 64'd3268106496, - 64'd143903696, 64'd99938729984, 64'd54692937728, - 64'd3410737920, - 64'd124915304, 64'd126815928320, 64'd52798849024, - 64'd3541361920, - 64'd106137392, 64'd152721162240, 64'd50806280192, - 64'd3659954688, - 64'd87605712, 64'd177607016448, 64'd48722604032, - 64'd3766520832, - 64'd69354872, 64'd201429811200, 64'd46555262976, - 64'd3861091584, - 64'd51418244, 64'd224149569536, 64'd44311724032, - 64'd3943725056, - 64'd33827940, 64'd245730066432, 64'd41999470592, - 64'd4014505728, - 64'd16614718, 64'd266138828800, 64'd39625990144, - 64'd4073542400, 64'd192039, 64'd285347086336, 64'd37198749696, - 64'd4120969216, 64'd16564378, 64'd303329837056, 64'd34725171200, - 64'd4156944384, 64'd32475822, 64'd320065765376, 64'd32212641792, - 64'd4181648384, 64'd47901400, 64'd335537209344, 64'd29668460544, - 64'd4195284480, 64'd62817684, 64'd349730144256, 64'd27099852800, - 64'd4198076672, 64'd77202808, 64'd362634149888, 64'd24513941504, - 64'd4190269952, 64'd91036512, 64'd374242344960, 64'd21917728768, - 64'd4172128256, 64'd104300136, 64'd384551321600, 64'd19318095872, - 64'd4143933952, 64'd116976656, 64'd393561014272, 64'd16721772544, - 64'd4105987072, 64'd129050688, 64'd401274732544, 64'd14135336960, - 64'd4058603776, 64'd140508480, 64'd407699062784, 64'd11565198336, - 64'd4002115584, 64'd151337968, 64'd412843671552, 64'd9017582592, - 64'd3936868608, 64'd161528704, 64'd416721371136, 64'd6498526720, - 64'd3863221248, 64'd171071872, 64'd419347922944, 64'd4013864704, - 64'd3781544960, 64'd179960336, 64'd420741906432, 64'd1569218048, - 64'd3692221952, 64'd188188528, 64'd420924719104, - 64'd830012288, - 64'd3595643392, 64'd195752544, 64'd419920347136, - 64'd3178654208, - 64'd3492210688, 64'd202650000, 64'd417755299840, - 64'd5471773184, - 64'd3382331648, 64'd208880144, 64'd414458576896, - 64'd7704678400, - 64'd3266421248, 64'd214443696, 64'd410061406208, - 64'd9872928768, - 64'd3144899584, 64'd219342912, 64'd404597145600, - 64'd11972338688, - 64'd3018191360, 64'd223581536, 64'd398101184512, - 64'd13998983168, - 64'd2886724096, 64'd227164720, 64'd390610878464, - 64'd15949202432, - 64'd2750928128, 64'd230099024, 64'd382165286912, - 64'd17819602944, - 64'd2611234560, 64'd232392368, 64'd372805107712, - 64'd19607060480, - 64'd2468074496, 64'd234054000, 64'd362572546048, - 64'd21308727296, - 64'd2321878272, 64'd235094384, 64'd351511117824, - 64'd22922024960, - 64'd2173074176, 64'd235525248, 64'd339665616896, - 64'd24444651520, - 64'd2022087680, 64'd235359472, 64'd327081918464, - 64'd25874577408, - 64'd1869340288, 64'd234611088, 64'd313806782464, - 64'd27210045440, - 64'd1715248896, 64'd233295104, 64'd299887853568, - 64'd28449574912, - 64'd1560224768, 64'd231427632, 64'd285373399040, - 64'd29591947264, - 64'd1404672512, 64'd229025680, 64'd270312259584, - 64'd30636220416, - 64'd1248989312, 64'd226107136, 64'd254753652736, - 64'd31581706240, - 64'd1093564416, 64'd222690768, 64'd238747090944, - 64'd32427984896, - 64'd938777984, 64'd218796064, 64'd222342234112, - 64'd33174886400, - 64'd785000704, 64'd214443280, 64'd205588758528, - 64'd33822494720, - 64'd632592832, 64'd209653280, 64'd188536242176, - 64'd34371137536, - 64'd481903776, 64'd204447520, 64'd171234033664, - 64'd34821386240, - 64'd333271232, 64'd198848016, 64'd153731137536, - 64'd35174043648, - 64'd187020832, 64'd192877200, 64'd136076091392, - 64'd35430129664, - 64'd43465508, 64'd186557968, 64'd118316892160, - 64'd35590901760, 64'd97094976, 64'd179913488, 64'd100500840448, - 64'd35657814016, 64'd234374464, 64'd172967280, 64'd82674450432, - 64'd35632529408, 64'd368100832, 64'd165743024, 64'd64883372032, - 64'd35516907520, 64'd498016320, 64'd158264592, 64'd47172263936, - 64'd35312996352, 64'd623877952, 64'd150555952, 64'd29584726016, - 64'd35023020032, 64'd745457600, 64'd142641120, 64'd12163198976, - 64'd34649366528, 64'd862542592, 64'd134544064, - 64'd5051114496, - 64'd34194597888, 64'd974935552, 64'd126288696, - 64'd22018322432, - 64'd33661411328, 64'd1082454656, 64'd117898832, - 64'd38699925504, - 64'd33052655616, 64'd1184934016, 64'd109398064, - 64'd55058870272, - 64'd32371302400, 64'd1282223232, 64'd100809776, - 64'd71059636224, - 64'd31620448256, 64'd1374188032, 64'd92157048, - 64'd86668263424, - 64'd30803302400, 64'd1460709888, 64'd83462640, - 64'd101852430336, - 64'd29923172352, 64'd1541685888, 64'd74748928, - 64'd116581498880, - 64'd28983453696, 64'd1617029120, 64'd66037868, - 64'd130826526720, - 64'd27987628032, 64'd1686668032, 64'd57350932, - 64'd144560357376, - 64'd26939242496, 64'd1750546944, 64'd48709088, - 64'd157757603840, - 64'd25841909760, 64'd1808625024, 64'd40132760, - 64'd170394714112, - 64'd24699285504, 64'd1860876672, 64'd31641770, - 64'd182449946624, - 64'd23515070464, 64'd1907291136, 64'd23255326, - 64'd193903460352, - 64'd22292994048, 64'd1947872512, 64'd14991971, - 64'd204737249280, - 64'd21036806144, 64'd1982638464, 64'd6869566, - 64'd214935207936, - 64'd19750268928, 64'd2011621248, - 64'd1094747, - 64'd224483082240, - 64'd18437144576, 64'd2034866304, - 64'd8884573, - 64'd233368535040, - 64'd17101187072, 64'd2052432256, - 64'd16484281, - 64'd241581080576, - 64'd15746132992, 64'd2064390784, - 64'd23879030, - 64'd249112100864, - 64'd14375695360, 64'd2070825600, - 64'd31054790, - 64'd255954829312, - 64'd12993552384, 64'd2071832192, - 64'd37998356, - 64'd262104301568, - 64'd11603337216, 64'd2067517952, - 64'd44697368, - 64'd267557404672, - 64'd10208634880, 64'd2058000640, - 64'd51140312, - 64'd272312778752, - 64'd8812969984, 64'd2043408768, - 64'd57316544, - 64'd276370784256, - 64'd7419803648, 64'd2023880448, - 64'd63216296, - 64'd279733567488, - 64'd6032520704, 64'd1999563520, - 64'd68830672, - 64'd282404847616, - 64'd4654428160, 64'd1970614144, - 64'd74151656, - 64'd284390031360, - 64'd3288744960, 64'd1937197184, - 64'd79172120, - 64'd285696163840, - 64'd1938598400, 64'd1899484800, - 64'd83885824, - 64'd286331731968, - 64'd607016704, 64'd1857656448, - 64'd88287392, - 64'd286306762752, 64'd703075968, 64'd1811898112, - 64'd92372336, - 64'd285632692224, 64'd1988864640, 64'd1762401536, - 64'd96137032, - 64'd284322398208, 64'd3247648256, 64'd1709363968, - 64'd99578704, - 64'd282389970944, 64'd4476844032, 64'd1652987392, - 64'd102695448, - 64'd279850876928, 64'd5673991680, 64'd1593477888, - 64'd105486176, - 64'd276721729536, 64'd6836756480, 64'd1531045248, - 64'd107950624, - 64'd273020223488, 64'd7962933760, 64'd1465902080, - 64'd110089344, - 64'd268765233152, 64'd9050448896, 64'd1398263424, - 64'd111903656, - 64'd263976550400, 64'd10097364992, 64'd1328346496, - 64'd113395672, - 64'd258674933760, 64'd11101879296, 64'd1256369408, - 64'd114568232, - 64'd252882010112, 64'd12062327808, 64'd1182551040, - 64'd115424912, - 64'd246620192768, 64'd12977186816, 64'd1107110656, - 64'd115969992, - 64'd239912648704, 64'd13845072896, 64'd1030267072, - 64'd116208416, - 64'd232783167488, 64'd14664743936, 64'd952238016, - 64'd116145800, - 64'd225256128512, 64'd15435101184, 64'd873240128, - 64'd115788360, - 64'd217356435456, 64'd16155185152, 64'd793487936, - 64'd115142944, - 64'd209109450752, 64'd16824177664, 64'd713193536, - 64'd114216936, - 64'd200540897280, 64'd17441402880, 64'd632566400, - 64'd113018280, - 64'd191676776448, 64'd18006323200, 64'd551812416, - 64'd111555416, - 64'd182543351808, 64'd18518538240, 64'd471133856, - 64'd109837272, - 64'd173167067136, 64'd18977785856, 64'd390728800, - 64'd107873208, - 64'd163574415360, 64'd19383932928, 64'd310790784, - 64'd105673032, - 64'd153791987712, 64'd19736985600, 64'd231508352, - 64'd103246896, - 64'd143846260736, 64'd20037074944, 64'd153064720, - 64'd100605320, - 64'd133763694592, 64'd20284461056, 64'd75637472, - 64'd97759152, - 64'd123570528256, 64'd20479520768, - 64'd601798, - 64'd94719512, - 64'd113292812288, 64'd20622761984, - 64'd75487776, - 64'd91497776, - 64'd102956302336, 64'd20714797056, - 64'd148861712, - 64'd88105536, - 64'd92586426368, 64'd20756363264, - 64'd220571664, - 64'd84554576, - 64'd82208210944, 64'd20748296192, - 64'd290472736, - 64'd80856832, - 64'd71846248448, 64'd20691544064, - 64'd358427360, - 64'd77024368, - 64'd61524611072, 64'd20587149312, - 64'd424305312, - 64'd73069320, - 64'd51266850816, 64'd20436252672, - 64'd487984128, - 64'd69003912, - 64'd41095909376, 64'd20240087040, - 64'd549349056, - 64'd64840380, - 64'd31034091520, 64'd19999971328, - 64'd608293248, - 64'd60590948, - 64'd21103032320, 64'd19717304320, - 64'd664717824, - 64'd56267824, - 64'd11323636736, 64'd19393564672, - 64'd718532160, - 64'd51883148, - 64'd1716058880, 64'd19030296576, - 64'd769653568, - 64'd47448976, 64'd7700338176, 64'd18629117952, - 64'd818007744, - 64'd42977236, 64'd16907015168, 64'd18191702016, - 64'd863528512, - 64'd38479724, 64'd25886285824, 64'd17719781376, - 64'd906157952, - 64'd33968056, 64'd34621337600, 64'd17215135744, - 64'd945846272, - 64'd29453662, 64'd43096268800, 64'd16679596032, - 64'd982551936, - 64'd24947746, 64'd51296092160, 64'd16115025920, - 64'd1016241344, - 64'd20461276, 64'd59206770688, 64'd15523328000, - 64'd1046889216, - 64'd16004951, 64'd66815217664, 64'd14906433536, - 64'd1074477824, - 64'd11589188, 64'd74109329408, 64'd14266298368, - 64'd1098997632, - 64'd7224101, 64'd81077968896, 64'd13604894720, - 64'd1120446464, - 64'd2919478, 64'd87711006720, 64'd12924210176, - 64'd1138829824, 64'd1315231, 64'd93999292416, 64'd12226242560, - 64'd1154160640, 64'd5470936, 64'd99934699520, 64'd11512990720, - 64'd1166458880, 64'd9538914, 64'd105510068224, 64'd10786453504, - 64'd1175751808, 64'd13510833, 64'd110719262720, 64'd10048623616, - 64'd1182073216, 64'd17378756, 64'd115557138432, 64'd9301481472, - 64'd1185463680, 64'd21135160, 64'd120019517440, 64'd8546993664, - 64'd1185970048, 64'd24772936, 64'd124103229440, 64'd7787105792, - 64'd1183645184, 64'd28285410, 64'd127806046208, 64'd7023740416, - 64'd1178548096, 64'd31666346, 64'd131126697984, 64'd6258790912, - 64'd1170743168, 64'd34909944, 64'd134064881664, 64'd5494117376, - 64'd1160300288, 64'd38010860, 64'd136621170688, 64'd4731544576, - 64'd1147294464, 64'd40964204, 64'd138797072384, 64'd3972856576, - 64'd1131805312, 64'd43765540, 64'd140594954240, 64'd3219794432, - 64'd1113917056, 64'd46410888, 64'd142018084864, 64'd2474051584, - 64'd1093718144, 64'd48896728, 64'd143070494720, 64'd1737271424, - 64'd1071300928, 64'd51220004, 64'd143757115392, 64'd1011044160, - 64'd1046761472, 64'd53378104, 64'd144083566592, 64'd296903744, - 64'd1020199040, 64'd55368892, 64'd144056270848, - 64'd403674336, - 64'd991715904, 64'd57190656, 64'd143682371584, - 64'd1089275904, - 64'd961417152, 64'd58842152, 64'd142969716736, - 64'd1758550016, - 64'd929410048, 64'd60322564, 64'd141926760448, - 64'd2410211328, - 64'd895804224, 64'd61631512, 64'd140562644992, - 64'd3043041536, - 64'd860710848, 64'd62769044, 64'd138887053312, - 64'd3655891456, - 64'd824242624, 64'd63735628, 64'd136910258176, - 64'd4247682048, - 64'd786513600, 64'd64532132, 64'd134643048448, - 64'd4817405952, - 64'd747638400, 64'd65159828, 64'd132096688128, - 64'd5364129280, - 64'd707732416, 64'd65620372, 64'd129282891776, - 64'd5886989824, - 64'd666911360, 64'd65915804, 64'd126213799936, - 64'd6385201664, - 64'd625290752, 64'd66048516, 64'd122901921792, - 64'd6858051584, - 64'd582985984, 64'd66021256, 64'd119360086016, - 64'd7304902656, - 64'd540111872, 64'd65837104, 64'd115601440768, - 64'd7725192704, - 64'd496782304, 64'd65499476, 64'd111639396352, - 64'd8118434304, - 64'd453110208, 64'd65012080, 64'd107487584256, - 64'd8484214272, - 64'd409207072, 64'd64378924, 64'd103159816192, - 64'd8822194176, - 64'd365182880, 64'd63604292, 64'd98670067712, - 64'd9132109824, - 64'd321145696, 64'd62692740, 64'd94032420864, - 64'd9413767168, - 64'd277201632, 64'd61649052, 64'd89261031424, - 64'd9667047424, - 64'd233454448, 64'd60478252, 64'd84370112512, - 64'd9891900416, - 64'd190005520, 64'd59185576, 64'd79373869056, - 64'd10088345600, - 64'd146953488, 64'd57776448, 64'd74286489600, - 64'd10256471040, - 64'd104394120, 64'd56256488, 64'd69122088960, - 64'd10396431360, - 64'd62420204, 64'd54631452, 64'd63894712320, - 64'd10508446720, - 64'd21121276, 64'd52907264, 64'd58618257408, - 64'd10592797696, 64'd19416466, 64'd51089960, 64'd53306470400, - 64'd10649829376, 64'd59110328, 64'd49185692};
	localparam logic signed[63:0] hb[0:1199] = {64'd4704787496960, 64'd4776038912, - 64'd6201745920, - 64'd12376386, 64'd4700013330432, 64'd14318410752, - 64'd6176088576, - 64'd37060376, 64'd4690473910272, 64'd23831724032, - 64'd6124879360, - 64'd61541484, 64'd4676189683712, 64'd33296730112, - 64'd6048317440, - 64'd85691840, 64'd4657188438016, 64'd42694332416, - 64'd5946690560, - 64'd109390016, 64'd4633509494784, 64'd52005650432, - 64'd5820371456, - 64'd132521128, 64'd4605200039936, 64'd61212069888, - 64'd5669813760, - 64'd154976880, 64'd4572317745152, 64'd70295289856, - 64'd5495548928, - 64'd176655632, 64'd4534928146432, 64'd79237382144, - 64'd5298182656, - 64'd197462448, 64'd4493106741248, 64'd88020836352, - 64'd5078390272, - 64'd217309056, 64'd4446936891392, 64'd96628596736, - 64'd4836913152, - 64'd236113952, 64'd4396510085120, 64'd105044131840, - 64'd4574555136, - 64'd253802304, 64'd4341927247872, 64'd113251434496, - 64'd4292176128, - 64'd270305984, 64'd4283295858688, 64'd121235111936, - 64'd3990691840, - 64'd285563488, 64'd4220731785216, 64'd128980369408, - 64'd3671066112, - 64'd299519904, 64'd4154357710848, 64'd136473083904, - 64'd3334309120, - 64'd312126848, 64'd4084303134720, 64'd143699820544, - 64'd2981470976, - 64'd323342368, 64'd4010704109568, 64'd150647848960, - 64'd2613640448, - 64'd333130880, 64'd3933703503872, 64'd157305192448, - 64'd2231937536, - 64'd341463008, 64'd3853449166848, 64'd163660644352, - 64'd1837512192, - 64'd348315488, 64'd3770094977024, 64'd169703784448, - 64'd1431538176, - 64'd353671104, 64'd3683799007232, 64'd175424978944, - 64'd1015210240, - 64'd357518464, 64'd3594725097472, 64'd180815462400, - 64'd589739520, - 64'd359851872, 64'd3503039971328, 64'd185867239424, - 64'd156349744, - 64'd360671232, 64'd3408915333120, 64'd190573232128, 64'd283726752, - 64'd359981728, 64'd3312525508608, 64'd194927149056, 64'd729252672, - 64'd357793824, 64'd3214047707136, 64'd198923616256, 64'd1178989696, - 64'd354122944, 64'd3113662283776, 64'd202558095360, 64'd1631701888, - 64'd348989408, 64'd3011550642176, 64'd205826899968, 64'd2086159488, - 64'd342418112, 64'd2907896545280, 64'd208727244800, 64'd2541142016, - 64'd334438336, 64'd2802885066752, 64'd211257163776, 64'd2995442432, - 64'd325083616, 64'd2696701280256, 64'd213415575552, 64'd3447869184, - 64'd314391488, 64'd2589531570176, 64'd215202234368, 64'd3897250048, - 64'd302403232, 64'd2481561010176, 64'd216617730048, 64'd4342434816, - 64'd289163680, 64'd2372975460352, 64'd217663455232, 64'd4782299136, - 64'd274721024, 64'd2263958683648, 64'd218341638144, 64'd5215745024, - 64'd259126464, 64'd2154694443008, 64'd218655309824, 64'd5641705984, - 64'd242434144, 64'd2045363617792, 64'd218608222208, 64'd6059147776, - 64'd224700832, 64'd1936145645568, 64'd218204946432, 64'd6467070976, - 64'd205985664, 64'd1827217211392, 64'd217450758144, 64'd6864514560, - 64'd186349936, 64'd1718752378880, 64'd216351637504, 64'd7250554880, - 64'd165856928, 64'd1610921934848, 64'd214914269184, 64'd7624310784, - 64'd144571552, 64'd1503893258240, 64'd213145993216, 64'd7984943616, - 64'd122560264, 64'd1397829795840, 64'd211054772224, 64'd8331659264, - 64'd99890704, 64'd1292890800128, 64'd208649191424, 64'd8663708672, - 64'd76631560, 64'd1189231460352, 64'd205938409472, 64'd8980389888, - 64'd52852316, 64'd1087001722880, 64'd202932142080, 64'd9281050624, - 64'd28623022, 64'd986346881024, 64'd199640612864, 64'd9565084672, - 64'd4014100, 64'd887406854144, 64'd196074520576, 64'd9831939072, 64'd20903884, 64'd790316253184, 64'd192245039104, 64'd10081110016, 64'd46060420, 64'd695203790848, 64'd188163735552, 64'd10312142848, 64'd71385240, 64'd602192478208, 64'd183842586624, 64'd10524638208, 64'd96808552, 64'd511399165952, 64'd179293913088, 64'd10718244864, 64'd122261184, 64'd422934413312, 64'd174530363392, 64'd10892664832, 64'd147674800, 64'd336902488064, 64'd169564848128, 64'd11047652352, 64'd172982048, 64'd253401055232, 64'd164410523648, 64'd11183011840, 64'd198116768, 64'd172521209856, 64'd159080792064, 64'd11298598912, 64'd223014128, 64'd94347255808, 64'd153589219328, 64'd11394321408, 64'd247610784, 64'd18956701696, 64'd147949502464, 64'd11470135296, 64'd271845024, - 64'd53579837440, 64'd142175469568, 64'd11526046720, 64'd295656928, - 64'd123198676992, 64'd136281006080, 64'd11562112000, 64'd318988480, - 64'd189843079168, 64'd130280062976, 64'd11578433536, 64'd341783712, - 64'd253463298048, 64'd124186583040, 64'd11575159808, 64'd363988800, - 64'd314016530432, 64'd118014500864, 64'd11552485376, 64'd385552160, - 64'd371466993664, 64'd111777677312, 64'd11510649856, 64'd406424608, - 64'd425785720832, 64'd105489899520, 64'd11449936896, 64'd426559392, - 64'd476950659072, 64'd99164839936, 64'd11370668032, 64'd445912288, - 64'd524946571264, 64'd92816015360, 64'd11273207808, 64'd464441728, - 64'd569764937728, 64'd86456786944, 64'd11157959680, 64'd482108768, - 64'd611403759616, 64'd80100278272, 64'd11025362944, 64'd498877216, - 64'd649867821056, 64'd73759424512, 64'd10875890688, 64'd514713696, - 64'd685167935488, 64'd67446861824, 64'd10710052864, 64'd529587616, - 64'd717321404416, 64'd61174980608, 64'd10528389120, 64'd543471232, - 64'd746351689728, 64'd54955843584, 64'd10331468800, 64'd556339776, - 64'd772288020480, 64'd48801189888, 64'd10119888896, 64'd568171200, - 64'd795165523968, 64'd42722418688, 64'd9894274048, 64'd578946624, - 64'd815024898048, 64'd36730548224, 64'd9655272448, 64'd588649792, - 64'd831912280064, 64'd30836209664, 64'd9403553792, 64'd597267584, - 64'd845879050240, 64'd25049632768, 64'd9139807232, 64'd604789568, - 64'd856981504000, 64'd19380617216, 64'd8864742400, 64'd611208448, - 64'd865280786432, 64'd13838529536, 64'd8579081728, 64'd616519488, - 64'd870842630144, 64'd8432279040, 64'd8283564544, 64'd620720832, - 64'd873737093120, 64'd3170313216, 64'd7978940416, 64'd623813568, - 64'd874038362112, - 64'd1939399552, 64'd7665970176, 64'd625801280, - 64'd871824359424, - 64'd6889375744, 64'd7345421312, 64'd626690240, - 64'd867176742912, - 64'd11672628224, 64'd7018067968, 64'd626489408, - 64'd860180578304, - 64'd16282670080, 64'd6684688384, 64'd625210304, - 64'd850923945984, - 64'd20713525248, 64'd6346062848, 64'd622866752, - 64'd839497809920, - 64'd24959727616, 64'd6002970624, 64'd619475072, - 64'd825995821056, - 64'd29016330240, 64'd5656191488, 64'd615053952, - 64'd810513793024, - 64'd32878905344, 64'd5306499072, 64'd609624128, - 64'd793149898752, - 64'd36543541248, 64'd4954663936, 64'd603208640, - 64'd774003818496, - 64'd40006840320, 64'd4601447424, 64'd595832512, - 64'd753177067520, - 64'd43265937408, 64'd4247603456, 64'd587522624, - 64'd730772340736, - 64'd46318465024, 64'd3893874944, 64'd578307904, - 64'd706893316096, - 64'd49162575872, 64'd3540992256, 64'd568218752, - 64'd681644720128, - 64'd51796918272, 64'd3189672704, 64'd557287488, - 64'd655131541504, - 64'd54220648448, 64'd2840618240, 64'd545547776, - 64'd627459227648, - 64'd56433414144, 64'd2494514432, 64'd533034752, - 64'd598733291520, - 64'd58435334144, 64'd2152028160, 64'd519784928, - 64'd569058918400, - 64'd60227010560, 64'd1813808128, 64'd505835904, - 64'd538541129728, - 64'd61809512448, 64'd1480481920, 64'd491226464, - 64'd507284029440, - 64'd63184347136, 64'd1152655872, 64'd475996352, - 64'd475391066112, - 64'd64353472512, 64'd830913536, 64'd460186112, - 64'd442964475904, - 64'd65319268352, 64'd515814912, 64'd443837152, - 64'd410105217024, - 64'd66084532224, 64'd207895440, 64'd426991392, - 64'd376912838656, - 64'd66652459008, - 64'd92334792, 64'd409691392, - 64'd343485054976, - 64'd67026620416, - 64'd384391904, 64'd391980032, - 64'd309917843456, - 64'd67210969088, - 64'd667818816, 64'd373900512, - 64'd276305018880, - 64'd67209797632, - 64'd942185920, 64'd355496224, - 64'd242738216960, - 64'd67027738624, - 64'd1207091584, 64'd336810688, - 64'd209306615808, - 64'd66669740032, - 64'd1462162688, 64'd317887360, - 64'd176096935936, - 64'd66141057024, - 64'd1707054720, 64'd298769568, - 64'd143193096192, - 64'd65447219200, - 64'd1941452544, 64'd279500384, - 64'd110676279296, - 64'd64594018304, - 64'd2165070336, 64'd260122560, - 64'd78624645120, - 64'd63587500032, - 64'd2377651712, 64'd240678480, - 64'd47113297920, - 64'd62433927168, - 64'd2578969600, 64'd221209920, - 64'd16214159360, - 64'd61139771392, - 64'd2768827136, 64'd201758064, 64'd14004141056, - 64'd59711692800, - 64'd2947056640, 64'd182363424, 64'd43476340736, - 64'd58156523520, - 64'd3113519360, 64'd163065696, 64'd72140636160, - 64'd56481234944, - 64'd3268106496, 64'd143903696, 64'd99938729984, - 64'd54692937728, - 64'd3410737920, 64'd124915304, 64'd126815928320, - 64'd52798849024, - 64'd3541361920, 64'd106137392, 64'd152721162240, - 64'd50806280192, - 64'd3659954688, 64'd87605712, 64'd177607016448, - 64'd48722604032, - 64'd3766520832, 64'd69354872, 64'd201429811200, - 64'd46555262976, - 64'd3861091584, 64'd51418244, 64'd224149569536, - 64'd44311724032, - 64'd3943725056, 64'd33827940, 64'd245730066432, - 64'd41999470592, - 64'd4014505728, 64'd16614718, 64'd266138828800, - 64'd39625990144, - 64'd4073542400, - 64'd192039, 64'd285347086336, - 64'd37198749696, - 64'd4120969216, - 64'd16564378, 64'd303329837056, - 64'd34725171200, - 64'd4156944384, - 64'd32475822, 64'd320065765376, - 64'd32212641792, - 64'd4181648384, - 64'd47901400, 64'd335537209344, - 64'd29668460544, - 64'd4195284480, - 64'd62817684, 64'd349730144256, - 64'd27099852800, - 64'd4198076672, - 64'd77202808, 64'd362634149888, - 64'd24513941504, - 64'd4190269952, - 64'd91036512, 64'd374242344960, - 64'd21917728768, - 64'd4172128256, - 64'd104300136, 64'd384551321600, - 64'd19318095872, - 64'd4143933952, - 64'd116976656, 64'd393561014272, - 64'd16721772544, - 64'd4105987072, - 64'd129050688, 64'd401274732544, - 64'd14135336960, - 64'd4058603776, - 64'd140508480, 64'd407699062784, - 64'd11565198336, - 64'd4002115584, - 64'd151337968, 64'd412843671552, - 64'd9017582592, - 64'd3936868608, - 64'd161528704, 64'd416721371136, - 64'd6498526720, - 64'd3863221248, - 64'd171071872, 64'd419347922944, - 64'd4013864704, - 64'd3781544960, - 64'd179960336, 64'd420741906432, - 64'd1569218048, - 64'd3692221952, - 64'd188188528, 64'd420924719104, 64'd830012288, - 64'd3595643392, - 64'd195752544, 64'd419920347136, 64'd3178654208, - 64'd3492210688, - 64'd202650000, 64'd417755299840, 64'd5471773184, - 64'd3382331648, - 64'd208880144, 64'd414458576896, 64'd7704678400, - 64'd3266421248, - 64'd214443696, 64'd410061406208, 64'd9872928768, - 64'd3144899584, - 64'd219342912, 64'd404597145600, 64'd11972338688, - 64'd3018191360, - 64'd223581536, 64'd398101184512, 64'd13998983168, - 64'd2886724096, - 64'd227164720, 64'd390610878464, 64'd15949202432, - 64'd2750928128, - 64'd230099024, 64'd382165286912, 64'd17819602944, - 64'd2611234560, - 64'd232392368, 64'd372805107712, 64'd19607060480, - 64'd2468074496, - 64'd234054000, 64'd362572546048, 64'd21308727296, - 64'd2321878272, - 64'd235094384, 64'd351511117824, 64'd22922024960, - 64'd2173074176, - 64'd235525248, 64'd339665616896, 64'd24444651520, - 64'd2022087680, - 64'd235359472, 64'd327081918464, 64'd25874577408, - 64'd1869340288, - 64'd234611088, 64'd313806782464, 64'd27210045440, - 64'd1715248896, - 64'd233295104, 64'd299887853568, 64'd28449574912, - 64'd1560224768, - 64'd231427632, 64'd285373399040, 64'd29591947264, - 64'd1404672512, - 64'd229025680, 64'd270312259584, 64'd30636220416, - 64'd1248989312, - 64'd226107136, 64'd254753652736, 64'd31581706240, - 64'd1093564416, - 64'd222690768, 64'd238747090944, 64'd32427984896, - 64'd938777984, - 64'd218796064, 64'd222342234112, 64'd33174886400, - 64'd785000704, - 64'd214443280, 64'd205588758528, 64'd33822494720, - 64'd632592832, - 64'd209653280, 64'd188536242176, 64'd34371137536, - 64'd481903776, - 64'd204447520, 64'd171234033664, 64'd34821386240, - 64'd333271232, - 64'd198848016, 64'd153731137536, 64'd35174043648, - 64'd187020832, - 64'd192877200, 64'd136076091392, 64'd35430129664, - 64'd43465508, - 64'd186557968, 64'd118316892160, 64'd35590901760, 64'd97094976, - 64'd179913488, 64'd100500840448, 64'd35657814016, 64'd234374464, - 64'd172967280, 64'd82674450432, 64'd35632529408, 64'd368100832, - 64'd165743024, 64'd64883372032, 64'd35516907520, 64'd498016320, - 64'd158264592, 64'd47172263936, 64'd35312996352, 64'd623877952, - 64'd150555952, 64'd29584726016, 64'd35023020032, 64'd745457600, - 64'd142641120, 64'd12163198976, 64'd34649366528, 64'd862542592, - 64'd134544064, - 64'd5051114496, 64'd34194597888, 64'd974935552, - 64'd126288696, - 64'd22018322432, 64'd33661411328, 64'd1082454656, - 64'd117898832, - 64'd38699925504, 64'd33052655616, 64'd1184934016, - 64'd109398064, - 64'd55058870272, 64'd32371302400, 64'd1282223232, - 64'd100809776, - 64'd71059636224, 64'd31620448256, 64'd1374188032, - 64'd92157048, - 64'd86668263424, 64'd30803302400, 64'd1460709888, - 64'd83462640, - 64'd101852430336, 64'd29923172352, 64'd1541685888, - 64'd74748928, - 64'd116581498880, 64'd28983453696, 64'd1617029120, - 64'd66037868, - 64'd130826526720, 64'd27987628032, 64'd1686668032, - 64'd57350932, - 64'd144560357376, 64'd26939242496, 64'd1750546944, - 64'd48709088, - 64'd157757603840, 64'd25841909760, 64'd1808625024, - 64'd40132760, - 64'd170394714112, 64'd24699285504, 64'd1860876672, - 64'd31641770, - 64'd182449946624, 64'd23515070464, 64'd1907291136, - 64'd23255326, - 64'd193903460352, 64'd22292994048, 64'd1947872512, - 64'd14991971, - 64'd204737249280, 64'd21036806144, 64'd1982638464, - 64'd6869566, - 64'd214935207936, 64'd19750268928, 64'd2011621248, 64'd1094747, - 64'd224483082240, 64'd18437144576, 64'd2034866304, 64'd8884573, - 64'd233368535040, 64'd17101187072, 64'd2052432256, 64'd16484281, - 64'd241581080576, 64'd15746132992, 64'd2064390784, 64'd23879030, - 64'd249112100864, 64'd14375695360, 64'd2070825600, 64'd31054790, - 64'd255954829312, 64'd12993552384, 64'd2071832192, 64'd37998356, - 64'd262104301568, 64'd11603337216, 64'd2067517952, 64'd44697368, - 64'd267557404672, 64'd10208634880, 64'd2058000640, 64'd51140312, - 64'd272312778752, 64'd8812969984, 64'd2043408768, 64'd57316544, - 64'd276370784256, 64'd7419803648, 64'd2023880448, 64'd63216296, - 64'd279733567488, 64'd6032520704, 64'd1999563520, 64'd68830672, - 64'd282404847616, 64'd4654428160, 64'd1970614144, 64'd74151656, - 64'd284390031360, 64'd3288744960, 64'd1937197184, 64'd79172120, - 64'd285696163840, 64'd1938598400, 64'd1899484800, 64'd83885824, - 64'd286331731968, 64'd607016704, 64'd1857656448, 64'd88287392, - 64'd286306762752, - 64'd703075968, 64'd1811898112, 64'd92372336, - 64'd285632692224, - 64'd1988864640, 64'd1762401536, 64'd96137032, - 64'd284322398208, - 64'd3247648256, 64'd1709363968, 64'd99578704, - 64'd282389970944, - 64'd4476844032, 64'd1652987392, 64'd102695448, - 64'd279850876928, - 64'd5673991680, 64'd1593477888, 64'd105486176, - 64'd276721729536, - 64'd6836756480, 64'd1531045248, 64'd107950624, - 64'd273020223488, - 64'd7962933760, 64'd1465902080, 64'd110089344, - 64'd268765233152, - 64'd9050448896, 64'd1398263424, 64'd111903656, - 64'd263976550400, - 64'd10097364992, 64'd1328346496, 64'd113395672, - 64'd258674933760, - 64'd11101879296, 64'd1256369408, 64'd114568232, - 64'd252882010112, - 64'd12062327808, 64'd1182551040, 64'd115424912, - 64'd246620192768, - 64'd12977186816, 64'd1107110656, 64'd115969992, - 64'd239912648704, - 64'd13845072896, 64'd1030267072, 64'd116208416, - 64'd232783167488, - 64'd14664743936, 64'd952238016, 64'd116145800, - 64'd225256128512, - 64'd15435101184, 64'd873240128, 64'd115788360, - 64'd217356435456, - 64'd16155185152, 64'd793487936, 64'd115142944, - 64'd209109450752, - 64'd16824177664, 64'd713193536, 64'd114216936, - 64'd200540897280, - 64'd17441402880, 64'd632566400, 64'd113018280, - 64'd191676776448, - 64'd18006323200, 64'd551812416, 64'd111555416, - 64'd182543351808, - 64'd18518538240, 64'd471133856, 64'd109837272, - 64'd173167067136, - 64'd18977785856, 64'd390728800, 64'd107873208, - 64'd163574415360, - 64'd19383932928, 64'd310790784, 64'd105673032, - 64'd153791987712, - 64'd19736985600, 64'd231508352, 64'd103246896, - 64'd143846260736, - 64'd20037074944, 64'd153064720, 64'd100605320, - 64'd133763694592, - 64'd20284461056, 64'd75637472, 64'd97759152, - 64'd123570528256, - 64'd20479520768, - 64'd601798, 64'd94719512, - 64'd113292812288, - 64'd20622761984, - 64'd75487776, 64'd91497776, - 64'd102956302336, - 64'd20714797056, - 64'd148861712, 64'd88105536, - 64'd92586426368, - 64'd20756363264, - 64'd220571664, 64'd84554576, - 64'd82208210944, - 64'd20748296192, - 64'd290472736, 64'd80856832, - 64'd71846248448, - 64'd20691544064, - 64'd358427360, 64'd77024368, - 64'd61524611072, - 64'd20587149312, - 64'd424305312, 64'd73069320, - 64'd51266850816, - 64'd20436252672, - 64'd487984128, 64'd69003912, - 64'd41095909376, - 64'd20240087040, - 64'd549349056, 64'd64840380, - 64'd31034091520, - 64'd19999971328, - 64'd608293248, 64'd60590948, - 64'd21103032320, - 64'd19717304320, - 64'd664717824, 64'd56267824, - 64'd11323636736, - 64'd19393564672, - 64'd718532160, 64'd51883148, - 64'd1716058880, - 64'd19030296576, - 64'd769653568, 64'd47448976, 64'd7700338176, - 64'd18629117952, - 64'd818007744, 64'd42977236, 64'd16907015168, - 64'd18191702016, - 64'd863528512, 64'd38479724, 64'd25886285824, - 64'd17719781376, - 64'd906157952, 64'd33968056, 64'd34621337600, - 64'd17215135744, - 64'd945846272, 64'd29453662, 64'd43096268800, - 64'd16679596032, - 64'd982551936, 64'd24947746, 64'd51296092160, - 64'd16115025920, - 64'd1016241344, 64'd20461276, 64'd59206770688, - 64'd15523328000, - 64'd1046889216, 64'd16004951, 64'd66815217664, - 64'd14906433536, - 64'd1074477824, 64'd11589188, 64'd74109329408, - 64'd14266298368, - 64'd1098997632, 64'd7224101, 64'd81077968896, - 64'd13604894720, - 64'd1120446464, 64'd2919478, 64'd87711006720, - 64'd12924210176, - 64'd1138829824, - 64'd1315231, 64'd93999292416, - 64'd12226242560, - 64'd1154160640, - 64'd5470936, 64'd99934699520, - 64'd11512990720, - 64'd1166458880, - 64'd9538914, 64'd105510068224, - 64'd10786453504, - 64'd1175751808, - 64'd13510833, 64'd110719262720, - 64'd10048623616, - 64'd1182073216, - 64'd17378756, 64'd115557138432, - 64'd9301481472, - 64'd1185463680, - 64'd21135160, 64'd120019517440, - 64'd8546993664, - 64'd1185970048, - 64'd24772936, 64'd124103229440, - 64'd7787105792, - 64'd1183645184, - 64'd28285410, 64'd127806046208, - 64'd7023740416, - 64'd1178548096, - 64'd31666346, 64'd131126697984, - 64'd6258790912, - 64'd1170743168, - 64'd34909944, 64'd134064881664, - 64'd5494117376, - 64'd1160300288, - 64'd38010860, 64'd136621170688, - 64'd4731544576, - 64'd1147294464, - 64'd40964204, 64'd138797072384, - 64'd3972856576, - 64'd1131805312, - 64'd43765540, 64'd140594954240, - 64'd3219794432, - 64'd1113917056, - 64'd46410888, 64'd142018084864, - 64'd2474051584, - 64'd1093718144, - 64'd48896728, 64'd143070494720, - 64'd1737271424, - 64'd1071300928, - 64'd51220004, 64'd143757115392, - 64'd1011044160, - 64'd1046761472, - 64'd53378104, 64'd144083566592, - 64'd296903744, - 64'd1020199040, - 64'd55368892, 64'd144056270848, 64'd403674336, - 64'd991715904, - 64'd57190656, 64'd143682371584, 64'd1089275904, - 64'd961417152, - 64'd58842152, 64'd142969716736, 64'd1758550016, - 64'd929410048, - 64'd60322564, 64'd141926760448, 64'd2410211328, - 64'd895804224, - 64'd61631512, 64'd140562644992, 64'd3043041536, - 64'd860710848, - 64'd62769044, 64'd138887053312, 64'd3655891456, - 64'd824242624, - 64'd63735628, 64'd136910258176, 64'd4247682048, - 64'd786513600, - 64'd64532132, 64'd134643048448, 64'd4817405952, - 64'd747638400, - 64'd65159828, 64'd132096688128, 64'd5364129280, - 64'd707732416, - 64'd65620372, 64'd129282891776, 64'd5886989824, - 64'd666911360, - 64'd65915804, 64'd126213799936, 64'd6385201664, - 64'd625290752, - 64'd66048516, 64'd122901921792, 64'd6858051584, - 64'd582985984, - 64'd66021256, 64'd119360086016, 64'd7304902656, - 64'd540111872, - 64'd65837104, 64'd115601440768, 64'd7725192704, - 64'd496782304, - 64'd65499476, 64'd111639396352, 64'd8118434304, - 64'd453110208, - 64'd65012080, 64'd107487584256, 64'd8484214272, - 64'd409207072, - 64'd64378924, 64'd103159816192, 64'd8822194176, - 64'd365182880, - 64'd63604292, 64'd98670067712, 64'd9132109824, - 64'd321145696, - 64'd62692740, 64'd94032420864, 64'd9413767168, - 64'd277201632, - 64'd61649052, 64'd89261031424, 64'd9667047424, - 64'd233454448, - 64'd60478252, 64'd84370112512, 64'd9891900416, - 64'd190005520, - 64'd59185576, 64'd79373869056, 64'd10088345600, - 64'd146953488, - 64'd57776448, 64'd74286489600, 64'd10256471040, - 64'd104394120, - 64'd56256488, 64'd69122088960, 64'd10396431360, - 64'd62420204, - 64'd54631452, 64'd63894712320, 64'd10508446720, - 64'd21121276, - 64'd52907264, 64'd58618257408, 64'd10592797696, 64'd19416466, - 64'd51089960, 64'd53306470400, 64'd10649829376, 64'd59110328, - 64'd49185692};
endpackage
`endif
