`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam N = 5;
	localparam M = 5;
	localparam real Lfr[0:4] = {0.9753731, 0.9753731, 0.95266646, 0.95266646, 0.9445697};
	localparam real Lfi[0:4] = {0.12202396, -0.12202396, 0.07174822, -0.07174822, 0.0};
	localparam real Lbr[0:4] = {0.9753731, 0.9753731, 0.95266646, 0.95266646, 0.9445697};
	localparam real Lbi[0:4] = {0.12202396, -0.12202396, 0.07174822, -0.07174822, 0.0};
	localparam real Wfr[0:4] = {-2.2506598e-05, -2.2506598e-05, -3.0707335e-05, -3.0707335e-05, -4.0910054e-05};
	localparam real Wfi[0:4] = {-7.40372e-05, 7.40372e-05, 3.5388293e-05, -3.5388293e-05, -0.0};
	localparam real Wbr[0:4] = {2.2506598e-05, 2.2506598e-05, 3.0707335e-05, 3.0707335e-05, 4.0910054e-05};
	localparam real Wbi[0:4] = {7.40372e-05, -7.40372e-05, -3.5388293e-05, 3.5388293e-05, 0.0};
	localparam real Ffr[0:4][0:124] = '{
		'{43.064934, -19.57931, -0.63658524, 0.6594977, -0.05817887, 33.13118, -20.100471, -0.14379226, 0.6291185, -0.06789542, 23.019352, -20.292555, 0.33459356, 0.5900158, -0.07623184, 12.8921585, -20.163696, 0.79164535, 0.54309005, -0.08310552, 2.907052, -19.726723, 1.2210006, 0.4893325, -0.08845934, -6.7860317, -18.998808, 1.6169409, 0.4298068, -0.09226163, -16.046743, -18.001055, 1.9744586, 0.3656301, -0.09450585, -24.74617, -16.758034, 2.2893105, 0.2979539, -0.095209815, -32.76845, -15.297284, 2.558058, 0.22794509, -0.094414614, -40.012135, -13.648795, 2.7780926, 0.1567673, -0.09218317, -46.391243, -11.844448, 2.9476495, 0.08556297, -0.088598564, -51.836117, -9.917465, 3.0658045, 0.015436394, -0.083762005, -56.29392, -7.9018493, 3.1324623, -0.05256209, -0.077790715, -59.72888, -5.831825, 3.148328, -0.1174506, -0.07081553, -62.122314, -3.7413075, 3.114871, -0.17832859, -0.06297843, -63.472282, -1.6633842, 3.034274, -0.23438805, -0.054429956, -63.79309, 0.3701702, 2.9093778, -0.28492293, -0.045326587, -63.114513, 2.3293407, 2.743613, -0.3293366, -0.035828132, -61.480797, 4.1862783, 2.5409281, -0.3671475, -0.026095117, -58.949505, 5.9156585, 2.3057103, -0.39799258, -0.016286282, -55.59016, 7.4949884, 2.042703, -0.42162895, -0.0065561924, -51.482777, 8.90486, 1.7569194, -0.4379337, 0.0029470313, -46.71625, 10.129144, 1.4535575, -0.44690174, 0.012083783, -41.386703, 11.155135, 1.1379114, -0.44864166, 0.020724846, -35.595726, 11.973628, 0.8152873, -0.44337055, 0.02875305},
		'{43.064934, -19.57931, -0.63658524, 0.6594977, -0.05817887, 33.13118, -20.100471, -0.14379226, 0.6291185, -0.06789542, 23.019352, -20.292555, 0.33459356, 0.5900158, -0.07623184, 12.8921585, -20.163696, 0.79164535, 0.54309005, -0.08310552, 2.907052, -19.726723, 1.2210006, 0.4893325, -0.08845934, -6.7860317, -18.998808, 1.6169409, 0.4298068, -0.09226163, -16.046743, -18.001055, 1.9744586, 0.3656301, -0.09450585, -24.74617, -16.758034, 2.2893105, 0.2979539, -0.095209815, -32.76845, -15.297284, 2.558058, 0.22794509, -0.094414614, -40.012135, -13.648795, 2.7780926, 0.1567673, -0.09218317, -46.391243, -11.844448, 2.9476495, 0.08556297, -0.088598564, -51.836117, -9.917465, 3.0658045, 0.015436394, -0.083762005, -56.29392, -7.9018493, 3.1324623, -0.05256209, -0.077790715, -59.72888, -5.831825, 3.148328, -0.1174506, -0.07081553, -62.122314, -3.7413075, 3.114871, -0.17832859, -0.06297843, -63.472282, -1.6633842, 3.034274, -0.23438805, -0.054429956, -63.79309, 0.3701702, 2.9093778, -0.28492293, -0.045326587, -63.114513, 2.3293407, 2.743613, -0.3293366, -0.035828132, -61.480797, 4.1862783, 2.5409281, -0.3671475, -0.026095117, -58.949505, 5.9156585, 2.3057103, -0.39799258, -0.016286282, -55.59016, 7.4949884, 2.042703, -0.42162895, -0.0065561924, -51.482777, 8.90486, 1.7569194, -0.4379337, 0.0029470313, -46.71625, 10.129144, 1.4535575, -0.44690174, 0.012083783, -41.386703, 11.155135, 1.1379114, -0.44864166, 0.020724846, -35.595726, 11.973628, 0.8152873, -0.44337055, 0.02875305},
		'{-192.66455, 36.105915, -3.934311, 0.2366365, 0.12143486, -174.71106, 35.66837, -4.1022806, 0.32208657, 0.09852771, -157.03372, 35.00548, -4.2252812, 0.39769903, 0.07689192, -139.73903, 34.14182, -4.3063293, 0.4637738, 0.05657638, -122.921364, 33.101288, -4.348487, 0.5206551, 0.037615955, -106.663345, 31.907013, -4.3548374, 0.56872517, 0.020032454, -91.036255, 30.581234, -4.328459, 0.60839784, 0.0038356187, -76.10048, 29.145226, -4.272403, 0.64011294, -0.010975915, -61.90603, 27.619217, -4.1896734, 0.6643306, -0.024413623, -48.493076, 26.022339, -4.0832105, 0.68152636, -0.036498126, -35.89251, 24.372574, -3.9558713, 0.69218594, -0.04725825, -24.12652, 22.686726, -3.810419, 0.6968011, -0.056730088, -13.209201, 20.980402, -3.6495094, 0.6958654, -0.0649561, -3.1471393, 19.267996, -3.4756804, 0.68987006, -0.07198424, 6.059969, 17.562689, -3.2913435, 0.679301, -0.07786713, 14.418718, 15.876462, -3.0987778, 0.6646356, -0.08266126, 21.941397, 14.220106, -2.9001245, 0.6463396, -0.08642625, 28.645395, 12.603253, -2.6973827, 0.6248652, -0.08922409, 34.552635, 11.034402, -2.4924068, 0.60064834, -0.09111853, 39.68902, 9.520952, -2.2869065, 0.57410735, -0.09217441, 44.083866, 8.069252, -2.0824456, 0.5456411, -0.09245713, 47.769432, 6.684636, -1.8804443, 0.5156281, -0.092032075, 50.780396, 5.37148, -1.68218, 0.48442498, -0.09096415, 53.153385, 4.133249, -1.4887918, 0.45236614, -0.08931738, 54.92655, 2.9725513, -1.3012825, 0.41976318, -0.087154426},
		'{-192.66455, 36.105915, -3.934311, 0.2366365, 0.12143486, -174.71106, 35.66837, -4.1022806, 0.32208657, 0.09852771, -157.03372, 35.00548, -4.2252812, 0.39769903, 0.07689192, -139.73903, 34.14182, -4.3063293, 0.4637738, 0.05657638, -122.921364, 33.101288, -4.348487, 0.5206551, 0.037615955, -106.663345, 31.907013, -4.3548374, 0.56872517, 0.020032454, -91.036255, 30.581234, -4.328459, 0.60839784, 0.0038356187, -76.10048, 29.145226, -4.272403, 0.64011294, -0.010975915, -61.90603, 27.619217, -4.1896734, 0.6643306, -0.024413623, -48.493076, 26.022339, -4.0832105, 0.68152636, -0.036498126, -35.89251, 24.372574, -3.9558713, 0.69218594, -0.04725825, -24.12652, 22.686726, -3.810419, 0.6968011, -0.056730088, -13.209201, 20.980402, -3.6495094, 0.6958654, -0.0649561, -3.1471393, 19.267996, -3.4756804, 0.68987006, -0.07198424, 6.059969, 17.562689, -3.2913435, 0.679301, -0.07786713, 14.418718, 15.876462, -3.0987778, 0.6646356, -0.08266126, 21.941397, 14.220106, -2.9001245, 0.6463396, -0.08642625, 28.645395, 12.603253, -2.6973827, 0.6248652, -0.08922409, 34.552635, 11.034402, -2.4924068, 0.60064834, -0.09111853, 39.68902, 9.520952, -2.2869065, 0.57410735, -0.09217441, 44.083866, 8.069252, -2.0824456, 0.5456411, -0.09245713, 47.769432, 6.684636, -1.8804443, 0.5156281, -0.092032075, 50.780396, 5.37148, -1.68218, 0.48442498, -0.09096415, 53.153385, 4.133249, -1.4887918, 0.45236614, -0.08931738, 54.92655, 2.9725513, -1.3012825, 0.41976318, -0.087154426},
		'{-297.21286, 33.897514, -8.959085, 1.6006142, -0.34366232, -280.73828, 32.018566, -8.462481, 1.5118917, -0.324613, -265.17688, 30.243767, -7.993403, 1.4280871, -0.3066196, -250.47804, 28.567347, -7.550327, 1.3489279, -0.28962362, -236.59398, 26.98385, -7.1318097, 1.2741565, -0.2735697, -223.4795, 25.488129, -6.7364917, 1.2035296, -0.25840566, -211.09196, 24.075314, -6.363086, 1.1368176, -0.24408215, -199.39108, 22.740812, -6.0103784, 1.0738035, -0.23055261, -188.33878, 21.480284, -5.6772213, 1.0142822, -0.21777302, -177.89911, 20.289625, -5.3625317, 0.9580603, -0.2057018, -168.03812, 19.164965, -5.0652847, 0.9049548, -0.1942997, -158.72371, 18.102646, -4.784515, 0.8547929, -0.1835296, -149.92561, 17.09921, -4.5193076, 0.80741143, -0.1733565, -141.61519, 16.151398, -4.268801, 0.7626564, -0.16374731, -133.76543, 15.256121, -4.0321803, 0.72038215, -0.15467075, -126.35077, 14.41047, -3.8086755, 0.68045115, -0.1460973, -119.347115, 13.611693, -3.5975595, 0.6427336, -0.13799909, -112.73167, 12.857193, -3.398146, 0.6071067, -0.13034977, -106.48292, 12.144516, -3.2097857, 0.57345456, -0.123124436, -100.58054, 11.471342, -3.0318663, 0.5416678, -0.116299614, -95.00533, 10.835482, -2.863809, 0.51164305, -0.1098531, -89.73916, 10.234868, -2.7050674, 0.4832825, -0.10376391, -84.76489, 9.667546, -2.5551248, 0.45649403, -0.098012246, -80.06635, 9.131672, -2.4134934, 0.43119043, -0.0925794, -75.62825, 8.625501, -2.279713, 0.40728945, -0.087447695}};
	localparam real Ffi[0:4][0:124] = '{
		'{72.71686, 8.222471, -3.910018, 0.11586089, 0.09136989, 76.181015, 5.6308327, -3.8914049, 0.19348212, 0.08202052, 78.34772, 3.0394237, -3.813118, 0.26548478, 0.07171574, 79.227165, 0.4883941, -3.6783843, 0.33094278, 0.060647495, 78.849205, -1.9840876, -3.4911973, 0.3890627, 0.04901307, 77.26212, -4.3423586, -3.2562287, 0.43919158, 0.037011873, 74.531334, -6.5537295, -2.9787323, 0.48082238, 0.024842255, 70.73778, -8.588892, -2.6644442, 0.5135969, 0.012698489, 65.9761, -10.4222555, -2.3194766, 0.5373061, 0.0007678861, 60.352776, -12.032224, -1.9502107, 0.5518887, -0.01077187, 53.984035, -13.401387, -1.5631891, 0.55742675, -0.02175515, 46.993732, -14.516659, -1.1650088, 0.5541398, -0.032030534, 39.511177, -15.369328, -0.7622167, 0.54237664, -0.041462693, 31.668932, -15.955044, -0.36121017, 0.5226058, -0.04993393, 23.60067, -16.273743, 0.031856783, 0.49540383, -0.057345405, 15.439047, -16.3295, 0.41116115, 0.46144322, -0.06361804, 7.3136916, -16.13033, 0.7712897, 0.42147836, -0.06869309, -0.6507079, -15.687919, 1.107309, 0.37633124, -0.07253232, -8.336166, -15.017339, 1.414826, 0.3268764, -0.07511797, -15.633002, -14.1366825, 1.6900374, 0.27402565, -0.07645228, -22.441263, -13.066688, 1.9297689, 0.21871263, -0.07655681, -28.671936, -11.830328, 2.1315033, 0.16187759, -0.07547147, -34.247967, -10.452377, 2.2933974, 0.10445263, -0.07325323, -39.10505, -8.95897, 2.414287, 0.04734757, -0.06997472, -43.192184, -7.3771443, 2.493683, -0.008563485, -0.06572253},
		'{-72.71686, -8.222471, 3.910018, -0.11586089, -0.09136989, -76.181015, -5.6308327, 3.8914049, -0.19348212, -0.08202052, -78.34772, -3.0394237, 3.813118, -0.26548478, -0.07171574, -79.227165, -0.4883941, 3.6783843, -0.33094278, -0.060647495, -78.849205, 1.9840876, 3.4911973, -0.3890627, -0.04901307, -77.26212, 4.3423586, 3.2562287, -0.43919158, -0.037011873, -74.531334, 6.5537295, 2.9787323, -0.48082238, -0.024842255, -70.73778, 8.588892, 2.6644442, -0.5135969, -0.012698489, -65.9761, 10.4222555, 2.3194766, -0.5373061, -0.0007678861, -60.352776, 12.032224, 1.9502107, -0.5518887, 0.01077187, -53.984035, 13.401387, 1.5631891, -0.55742675, 0.02175515, -46.993732, 14.516659, 1.1650088, -0.5541398, 0.032030534, -39.511177, 15.369328, 0.7622167, -0.54237664, 0.041462693, -31.668932, 15.955044, 0.36121017, -0.5226058, 0.04993393, -23.60067, 16.273743, -0.031856783, -0.49540383, 0.057345405, -15.439047, 16.3295, -0.41116115, -0.46144322, 0.06361804, -7.3136916, 16.13033, -0.7712897, -0.42147836, 0.06869309, 0.6507079, 15.687919, -1.107309, -0.37633124, 0.07253232, 8.336166, 15.017339, -1.414826, -0.3268764, 0.07511797, 15.633002, 14.1366825, -1.6900374, -0.27402565, 0.07645228, 22.441263, 13.066688, -1.9297689, -0.21871263, 0.07655681, 28.671936, 11.830328, -2.1315033, -0.16187759, 0.07547147, 34.247967, 10.452377, -2.2933974, -0.10445263, 0.07325323, 39.10505, 8.95897, -2.414287, -0.04734757, 0.06997472, 43.192184, 7.3771443, -2.493683, 0.008563485, 0.06572253},
		'{-123.12489, -17.721321, 4.936633, -1.3470846, 0.2391586, -131.12029, -14.291972, 4.420685, -1.2663441, 0.23655112, -137.44911, -11.05634, 3.9171069, -1.1832944, 0.2324235, -142.21004, -8.021423, 3.42854, -1.0987507, 0.22693892, -145.50476, -5.192126, 2.9572835, -1.0134679, 0.22025634, -147.43689, -2.5714054, 2.5053084, -0.9281408, 0.2125297, -148.11108, -0.16042013, 2.0742714, -0.8434036, 0.20390722, -147.63216, 2.0413222, 1.6655296, -0.75983083, 0.19453076, -146.10426, 4.035817, 1.2801569, -0.67793834, 0.18453543, -143.63028, 5.8264174, 0.9189608, -0.5981846, 0.17404906, -140.31104, 7.417689, 0.58250004, -0.5209721, 0.16319203, -136.24484, 8.815272, 0.2711015, -0.4466495, 0.15207689, -131.52692, 10.025746, -0.015121497, -0.37551373, 0.14080825, -126.24902, 11.056499, -0.27625155, -0.30781224, 0.12948282, -120.49901, 11.9156, -0.51254946, -0.24374545, 0.11818919, -114.36057, 12.611684, -0.7244367, -0.18346946, 0.10700805, -107.91296, 13.153835, -0.9124783, -0.12709878, 0.096012175, -101.2308, 13.551485, -1.0773662, -0.07470902, 0.08526665, -94.38393, 13.814306, -1.2199031, -0.026339812, 0.074829005, -87.43731, 13.952125, -1.3409865, 0.018002395, 0.06474949, -80.45097, 13.974832, -1.4415944, 0.058341455, 0.055071317, -73.48, 13.892308, -1.5227703, 0.09472873, 0.04583096, -66.57456, 13.714346, -1.5856107, 0.12724029, 0.03705848, -59.77995, 13.450592, -1.6312516, 0.15597418, 0.028777855, -53.13669, 13.11048, -1.6608567, 0.18104783, 0.021007333},
		'{123.12489, 17.721321, -4.936633, 1.3470846, -0.2391586, 131.12029, 14.291972, -4.420685, 1.2663441, -0.23655112, 137.44911, 11.05634, -3.9171069, 1.1832944, -0.2324235, 142.21004, 8.021423, -3.42854, 1.0987507, -0.22693892, 145.50476, 5.192126, -2.9572835, 1.0134679, -0.22025634, 147.43689, 2.5714054, -2.5053084, 0.9281408, -0.2125297, 148.11108, 0.16042013, -2.0742714, 0.8434036, -0.20390722, 147.63216, -2.0413222, -1.6655296, 0.75983083, -0.19453076, 146.10426, -4.035817, -1.2801569, 0.67793834, -0.18453543, 143.63028, -5.8264174, -0.9189608, 0.5981846, -0.17404906, 140.31104, -7.417689, -0.58250004, 0.5209721, -0.16319203, 136.24484, -8.815272, -0.2711015, 0.4466495, -0.15207689, 131.52692, -10.025746, 0.015121497, 0.37551373, -0.14080825, 126.24902, -11.056499, 0.27625155, 0.30781224, -0.12948282, 120.49901, -11.9156, 0.51254946, 0.24374545, -0.11818919, 114.36057, -12.611684, 0.7244367, 0.18346946, -0.10700805, 107.91296, -13.153835, 0.9124783, 0.12709878, -0.096012175, 101.2308, -13.551485, 1.0773662, 0.07470902, -0.08526665, 94.38393, -13.814306, 1.2199031, 0.026339812, -0.074829005, 87.43731, -13.952125, 1.3409865, -0.018002395, -0.06474949, 80.45097, -13.974832, 1.4415944, -0.058341455, -0.055071317, 73.48, -13.892308, 1.5227703, -0.09472873, -0.04583096, 66.57456, -13.714346, 1.5856107, -0.12724029, -0.03705848, 59.77995, -13.450592, 1.6312516, -0.15597418, -0.028777855, 53.13669, -13.11048, 1.6608567, -0.18104783, -0.021007333},
		'{1.5015588e-11, 2.1104364e-12, -7.663234e-13, 6.098396e-14, 3.869166e-15, 1.418327e-11, 1.9934542e-12, -7.238459e-13, 5.76036e-14, 3.654697e-15, 1.3397087e-11, 1.8829565e-12, -6.8372294e-13, 5.4410615e-14, 3.452116e-15, 1.26544825e-11, 1.7785837e-12, -6.45824e-13, 5.1394622e-14, 3.2607643e-15, 1.1953041e-11, 1.6799963e-12, -6.1002576e-13, 4.8545803e-14, 3.0800191e-15, 1.1290481e-11, 1.5868736e-12, -5.762119e-13, 4.5854894e-14, 2.9092928e-15, 1.0664646e-11, 1.4989128e-12, -5.442723e-13, 4.3313145e-14, 2.74803e-15, 1.0073502e-11, 1.4158276e-12, -5.1410314e-13, 4.0912284e-14, 2.5957058e-15, 9.515125e-12, 1.3373479e-12, -4.8560624e-13, 3.8644506e-14, 2.4518252e-15, 8.987699e-12, 1.2632184e-12, -4.5868897e-13, 3.650243e-14, 2.3159198e-15, 8.489509e-12, 1.1931978e-12, -4.332637e-13, 3.447909e-14, 2.1875477e-15, 8.018933e-12, 1.1270585e-12, -4.0924778e-13, 3.2567905e-14, 2.0662913e-15, 7.574441e-12, 1.0645854e-12, -3.8656304e-13, 3.0762658e-14, 1.9517562e-15, 7.1545873e-12, 1.0055751e-12, -3.6513576e-13, 2.9057475e-14, 1.8435698e-15, 6.7580065e-12, 9.498358e-13, -3.4489618e-13, 2.744681e-14, 1.7413803e-15, 6.3834086e-12, 8.971861e-13, -3.257785e-13, 2.5925425e-14, 1.6448551e-15, 6.0295744e-12, 8.474548e-13, -3.0772048e-13, 2.4488373e-14, 1.5536802e-15, 5.6953535e-12, 8.004802e-13, -2.9066346e-13, 2.3130976e-14, 1.4675593e-15, 5.379658e-12, 7.561093e-13, -2.745519e-13, 2.1848818e-14, 1.3862121e-15, 5.081462e-12, 7.1419796e-13, -2.593334e-13, 2.0637732e-14, 1.309374e-15, 4.7997955e-12, 6.746098e-13, -2.4495849e-13, 1.9493777e-14, 1.236795e-15, 4.5337414e-12, 6.37216e-13, -2.3138037e-13, 1.841323e-14, 1.1682392e-15, 4.282435e-12, 6.018949e-13, -2.185549e-13, 1.7392582e-14, 1.1034833e-15, 4.045058e-12, 5.685317e-13, -2.0644033e-13, 1.6428506e-14, 1.0423169e-15, 3.8208395e-12, 5.3701786e-13, -1.9499728e-13, 1.5517869e-14, 9.84541e-16}};
	localparam real Fbr[0:4][0:124] = '{
		'{-43.064934, -19.57931, 0.63658524, 0.6594977, 0.05817887, -33.13118, -20.100471, 0.14379226, 0.6291185, 0.06789542, -23.019352, -20.292555, -0.33459356, 0.5900158, 0.07623184, -12.8921585, -20.163696, -0.79164535, 0.54309005, 0.08310552, -2.907052, -19.726723, -1.2210006, 0.4893325, 0.08845934, 6.7860317, -18.998808, -1.6169409, 0.4298068, 0.09226163, 16.046743, -18.001055, -1.9744586, 0.3656301, 0.09450585, 24.74617, -16.758034, -2.2893105, 0.2979539, 0.095209815, 32.76845, -15.297284, -2.558058, 0.22794509, 0.094414614, 40.012135, -13.648795, -2.7780926, 0.1567673, 0.09218317, 46.391243, -11.844448, -2.9476495, 0.08556297, 0.088598564, 51.836117, -9.917465, -3.0658045, 0.015436394, 0.083762005, 56.29392, -7.9018493, -3.1324623, -0.05256209, 0.077790715, 59.72888, -5.831825, -3.148328, -0.1174506, 0.07081553, 62.122314, -3.7413075, -3.114871, -0.17832859, 0.06297843, 63.472282, -1.6633842, -3.034274, -0.23438805, 0.054429956, 63.79309, 0.3701702, -2.9093778, -0.28492293, 0.045326587, 63.114513, 2.3293407, -2.743613, -0.3293366, 0.035828132, 61.480797, 4.1862783, -2.5409281, -0.3671475, 0.026095117, 58.949505, 5.9156585, -2.3057103, -0.39799258, 0.016286282, 55.59016, 7.4949884, -2.042703, -0.42162895, 0.0065561924, 51.482777, 8.90486, -1.7569194, -0.4379337, -0.0029470313, 46.71625, 10.129144, -1.4535575, -0.44690174, -0.012083783, 41.386703, 11.155135, -1.1379114, -0.44864166, -0.020724846, 35.595726, 11.973628, -0.8152873, -0.44337055, -0.02875305},
		'{-43.064934, -19.57931, 0.63658524, 0.6594977, 0.05817887, -33.13118, -20.100471, 0.14379226, 0.6291185, 0.06789542, -23.019352, -20.292555, -0.33459356, 0.5900158, 0.07623184, -12.8921585, -20.163696, -0.79164535, 0.54309005, 0.08310552, -2.907052, -19.726723, -1.2210006, 0.4893325, 0.08845934, 6.7860317, -18.998808, -1.6169409, 0.4298068, 0.09226163, 16.046743, -18.001055, -1.9744586, 0.3656301, 0.09450585, 24.74617, -16.758034, -2.2893105, 0.2979539, 0.095209815, 32.76845, -15.297284, -2.558058, 0.22794509, 0.094414614, 40.012135, -13.648795, -2.7780926, 0.1567673, 0.09218317, 46.391243, -11.844448, -2.9476495, 0.08556297, 0.088598564, 51.836117, -9.917465, -3.0658045, 0.015436394, 0.083762005, 56.29392, -7.9018493, -3.1324623, -0.05256209, 0.077790715, 59.72888, -5.831825, -3.148328, -0.1174506, 0.07081553, 62.122314, -3.7413075, -3.114871, -0.17832859, 0.06297843, 63.472282, -1.6633842, -3.034274, -0.23438805, 0.054429956, 63.79309, 0.3701702, -2.9093778, -0.28492293, 0.045326587, 63.114513, 2.3293407, -2.743613, -0.3293366, 0.035828132, 61.480797, 4.1862783, -2.5409281, -0.3671475, 0.026095117, 58.949505, 5.9156585, -2.3057103, -0.39799258, 0.016286282, 55.59016, 7.4949884, -2.042703, -0.42162895, 0.0065561924, 51.482777, 8.90486, -1.7569194, -0.4379337, -0.0029470313, 46.71625, 10.129144, -1.4535575, -0.44690174, -0.012083783, 41.386703, 11.155135, -1.1379114, -0.44864166, -0.020724846, 35.595726, 11.973628, -0.8152873, -0.44337055, -0.02875305},
		'{192.66455, 36.105915, 3.934311, 0.2366365, -0.12143486, 174.71106, 35.66837, 4.1022806, 0.32208657, -0.09852771, 157.03372, 35.00548, 4.2252812, 0.39769903, -0.07689192, 139.73903, 34.14182, 4.3063293, 0.4637738, -0.05657638, 122.921364, 33.101288, 4.348487, 0.5206551, -0.037615955, 106.663345, 31.907013, 4.3548374, 0.56872517, -0.020032454, 91.036255, 30.581234, 4.328459, 0.60839784, -0.0038356187, 76.10048, 29.145226, 4.272403, 0.64011294, 0.010975915, 61.90603, 27.619217, 4.1896734, 0.6643306, 0.024413623, 48.493076, 26.022339, 4.0832105, 0.68152636, 0.036498126, 35.89251, 24.372574, 3.9558713, 0.69218594, 0.04725825, 24.12652, 22.686726, 3.810419, 0.6968011, 0.056730088, 13.209201, 20.980402, 3.6495094, 0.6958654, 0.0649561, 3.1471393, 19.267996, 3.4756804, 0.68987006, 0.07198424, -6.059969, 17.562689, 3.2913435, 0.679301, 0.07786713, -14.418718, 15.876462, 3.0987778, 0.6646356, 0.08266126, -21.941397, 14.220106, 2.9001245, 0.6463396, 0.08642625, -28.645395, 12.603253, 2.6973827, 0.6248652, 0.08922409, -34.552635, 11.034402, 2.4924068, 0.60064834, 0.09111853, -39.68902, 9.520952, 2.2869065, 0.57410735, 0.09217441, -44.083866, 8.069252, 2.0824456, 0.5456411, 0.09245713, -47.769432, 6.684636, 1.8804443, 0.5156281, 0.092032075, -50.780396, 5.37148, 1.68218, 0.48442498, 0.09096415, -53.153385, 4.133249, 1.4887918, 0.45236614, 0.08931738, -54.92655, 2.9725513, 1.3012825, 0.41976318, 0.087154426},
		'{192.66455, 36.105915, 3.934311, 0.2366365, -0.12143486, 174.71106, 35.66837, 4.1022806, 0.32208657, -0.09852771, 157.03372, 35.00548, 4.2252812, 0.39769903, -0.07689192, 139.73903, 34.14182, 4.3063293, 0.4637738, -0.05657638, 122.921364, 33.101288, 4.348487, 0.5206551, -0.037615955, 106.663345, 31.907013, 4.3548374, 0.56872517, -0.020032454, 91.036255, 30.581234, 4.328459, 0.60839784, -0.0038356187, 76.10048, 29.145226, 4.272403, 0.64011294, 0.010975915, 61.90603, 27.619217, 4.1896734, 0.6643306, 0.024413623, 48.493076, 26.022339, 4.0832105, 0.68152636, 0.036498126, 35.89251, 24.372574, 3.9558713, 0.69218594, 0.04725825, 24.12652, 22.686726, 3.810419, 0.6968011, 0.056730088, 13.209201, 20.980402, 3.6495094, 0.6958654, 0.0649561, 3.1471393, 19.267996, 3.4756804, 0.68987006, 0.07198424, -6.059969, 17.562689, 3.2913435, 0.679301, 0.07786713, -14.418718, 15.876462, 3.0987778, 0.6646356, 0.08266126, -21.941397, 14.220106, 2.9001245, 0.6463396, 0.08642625, -28.645395, 12.603253, 2.6973827, 0.6248652, 0.08922409, -34.552635, 11.034402, 2.4924068, 0.60064834, 0.09111853, -39.68902, 9.520952, 2.2869065, 0.57410735, 0.09217441, -44.083866, 8.069252, 2.0824456, 0.5456411, 0.09245713, -47.769432, 6.684636, 1.8804443, 0.5156281, 0.092032075, -50.780396, 5.37148, 1.68218, 0.48442498, 0.09096415, -53.153385, 4.133249, 1.4887918, 0.45236614, 0.08931738, -54.92655, 2.9725513, 1.3012825, 0.41976318, 0.087154426},
		'{297.21286, 33.897514, 8.959085, 1.6006142, 0.34366232, 280.73828, 32.018566, 8.462481, 1.5118917, 0.324613, 265.17688, 30.243767, 7.993403, 1.4280871, 0.3066196, 250.47804, 28.567347, 7.550327, 1.3489279, 0.28962362, 236.59398, 26.98385, 7.1318097, 1.2741565, 0.2735697, 223.4795, 25.488129, 6.7364917, 1.2035296, 0.25840566, 211.09196, 24.075314, 6.363086, 1.1368176, 0.24408215, 199.39108, 22.740812, 6.0103784, 1.0738035, 0.23055261, 188.33878, 21.480284, 5.6772213, 1.0142822, 0.21777302, 177.89911, 20.289625, 5.3625317, 0.9580603, 0.2057018, 168.03812, 19.164965, 5.0652847, 0.9049548, 0.1942997, 158.72371, 18.102646, 4.784515, 0.8547929, 0.1835296, 149.92561, 17.09921, 4.5193076, 0.80741143, 0.1733565, 141.61519, 16.151398, 4.268801, 0.7626564, 0.16374731, 133.76543, 15.256121, 4.0321803, 0.72038215, 0.15467075, 126.35077, 14.41047, 3.8086755, 0.68045115, 0.1460973, 119.347115, 13.611693, 3.5975595, 0.6427336, 0.13799909, 112.73167, 12.857193, 3.398146, 0.6071067, 0.13034977, 106.48292, 12.144516, 3.2097857, 0.57345456, 0.123124436, 100.58054, 11.471342, 3.0318663, 0.5416678, 0.116299614, 95.00533, 10.835482, 2.863809, 0.51164305, 0.1098531, 89.73916, 10.234868, 2.7050674, 0.4832825, 0.10376391, 84.76489, 9.667546, 2.5551248, 0.45649403, 0.098012246, 80.06635, 9.131672, 2.4134934, 0.43119043, 0.0925794, 75.62825, 8.625501, 2.279713, 0.40728945, 0.087447695}};
	localparam real Fbi[0:4][0:124] = '{
		'{-72.71686, 8.222471, 3.910018, 0.11586089, -0.09136989, -76.181015, 5.6308327, 3.8914049, 0.19348212, -0.08202052, -78.34772, 3.0394237, 3.813118, 0.26548478, -0.07171574, -79.227165, 0.4883941, 3.6783843, 0.33094278, -0.060647495, -78.849205, -1.9840876, 3.4911973, 0.3890627, -0.04901307, -77.26212, -4.3423586, 3.2562287, 0.43919158, -0.037011873, -74.531334, -6.5537295, 2.9787323, 0.48082238, -0.024842255, -70.73778, -8.588892, 2.6644442, 0.5135969, -0.012698489, -65.9761, -10.4222555, 2.3194766, 0.5373061, -0.0007678861, -60.352776, -12.032224, 1.9502107, 0.5518887, 0.01077187, -53.984035, -13.401387, 1.5631891, 0.55742675, 0.02175515, -46.993732, -14.516659, 1.1650088, 0.5541398, 0.032030534, -39.511177, -15.369328, 0.7622167, 0.54237664, 0.041462693, -31.668932, -15.955044, 0.36121017, 0.5226058, 0.04993393, -23.60067, -16.273743, -0.031856783, 0.49540383, 0.057345405, -15.439047, -16.3295, -0.41116115, 0.46144322, 0.06361804, -7.3136916, -16.13033, -0.7712897, 0.42147836, 0.06869309, 0.6507079, -15.687919, -1.107309, 0.37633124, 0.07253232, 8.336166, -15.017339, -1.414826, 0.3268764, 0.07511797, 15.633002, -14.1366825, -1.6900374, 0.27402565, 0.07645228, 22.441263, -13.066688, -1.9297689, 0.21871263, 0.07655681, 28.671936, -11.830328, -2.1315033, 0.16187759, 0.07547147, 34.247967, -10.452377, -2.2933974, 0.10445263, 0.07325323, 39.10505, -8.95897, -2.414287, 0.04734757, 0.06997472, 43.192184, -7.3771443, -2.493683, -0.008563485, 0.06572253},
		'{72.71686, -8.222471, -3.910018, -0.11586089, 0.09136989, 76.181015, -5.6308327, -3.8914049, -0.19348212, 0.08202052, 78.34772, -3.0394237, -3.813118, -0.26548478, 0.07171574, 79.227165, -0.4883941, -3.6783843, -0.33094278, 0.060647495, 78.849205, 1.9840876, -3.4911973, -0.3890627, 0.04901307, 77.26212, 4.3423586, -3.2562287, -0.43919158, 0.037011873, 74.531334, 6.5537295, -2.9787323, -0.48082238, 0.024842255, 70.73778, 8.588892, -2.6644442, -0.5135969, 0.012698489, 65.9761, 10.4222555, -2.3194766, -0.5373061, 0.0007678861, 60.352776, 12.032224, -1.9502107, -0.5518887, -0.01077187, 53.984035, 13.401387, -1.5631891, -0.55742675, -0.02175515, 46.993732, 14.516659, -1.1650088, -0.5541398, -0.032030534, 39.511177, 15.369328, -0.7622167, -0.54237664, -0.041462693, 31.668932, 15.955044, -0.36121017, -0.5226058, -0.04993393, 23.60067, 16.273743, 0.031856783, -0.49540383, -0.057345405, 15.439047, 16.3295, 0.41116115, -0.46144322, -0.06361804, 7.3136916, 16.13033, 0.7712897, -0.42147836, -0.06869309, -0.6507079, 15.687919, 1.107309, -0.37633124, -0.07253232, -8.336166, 15.017339, 1.414826, -0.3268764, -0.07511797, -15.633002, 14.1366825, 1.6900374, -0.27402565, -0.07645228, -22.441263, 13.066688, 1.9297689, -0.21871263, -0.07655681, -28.671936, 11.830328, 2.1315033, -0.16187759, -0.07547147, -34.247967, 10.452377, 2.2933974, -0.10445263, -0.07325323, -39.10505, 8.95897, 2.414287, -0.04734757, -0.06997472, -43.192184, 7.3771443, 2.493683, 0.008563485, -0.06572253},
		'{123.12489, -17.721321, -4.936633, -1.3470846, -0.2391586, 131.12029, -14.291972, -4.420685, -1.2663441, -0.23655112, 137.44911, -11.05634, -3.9171069, -1.1832944, -0.2324235, 142.21004, -8.021423, -3.42854, -1.0987507, -0.22693892, 145.50476, -5.192126, -2.9572835, -1.0134679, -0.22025634, 147.43689, -2.5714054, -2.5053084, -0.9281408, -0.2125297, 148.11108, -0.16042013, -2.0742714, -0.8434036, -0.20390722, 147.63216, 2.0413222, -1.6655296, -0.75983083, -0.19453076, 146.10426, 4.035817, -1.2801569, -0.67793834, -0.18453543, 143.63028, 5.8264174, -0.9189608, -0.5981846, -0.17404906, 140.31104, 7.417689, -0.58250004, -0.5209721, -0.16319203, 136.24484, 8.815272, -0.2711015, -0.4466495, -0.15207689, 131.52692, 10.025746, 0.015121497, -0.37551373, -0.14080825, 126.24902, 11.056499, 0.27625155, -0.30781224, -0.12948282, 120.49901, 11.9156, 0.51254946, -0.24374545, -0.11818919, 114.36057, 12.611684, 0.7244367, -0.18346946, -0.10700805, 107.91296, 13.153835, 0.9124783, -0.12709878, -0.096012175, 101.2308, 13.551485, 1.0773662, -0.07470902, -0.08526665, 94.38393, 13.814306, 1.2199031, -0.026339812, -0.074829005, 87.43731, 13.952125, 1.3409865, 0.018002395, -0.06474949, 80.45097, 13.974832, 1.4415944, 0.058341455, -0.055071317, 73.48, 13.892308, 1.5227703, 0.09472873, -0.04583096, 66.57456, 13.714346, 1.5856107, 0.12724029, -0.03705848, 59.77995, 13.450592, 1.6312516, 0.15597418, -0.028777855, 53.13669, 13.11048, 1.6608567, 0.18104783, -0.021007333},
		'{-123.12489, 17.721321, 4.936633, 1.3470846, 0.2391586, -131.12029, 14.291972, 4.420685, 1.2663441, 0.23655112, -137.44911, 11.05634, 3.9171069, 1.1832944, 0.2324235, -142.21004, 8.021423, 3.42854, 1.0987507, 0.22693892, -145.50476, 5.192126, 2.9572835, 1.0134679, 0.22025634, -147.43689, 2.5714054, 2.5053084, 0.9281408, 0.2125297, -148.11108, 0.16042013, 2.0742714, 0.8434036, 0.20390722, -147.63216, -2.0413222, 1.6655296, 0.75983083, 0.19453076, -146.10426, -4.035817, 1.2801569, 0.67793834, 0.18453543, -143.63028, -5.8264174, 0.9189608, 0.5981846, 0.17404906, -140.31104, -7.417689, 0.58250004, 0.5209721, 0.16319203, -136.24484, -8.815272, 0.2711015, 0.4466495, 0.15207689, -131.52692, -10.025746, -0.015121497, 0.37551373, 0.14080825, -126.24902, -11.056499, -0.27625155, 0.30781224, 0.12948282, -120.49901, -11.9156, -0.51254946, 0.24374545, 0.11818919, -114.36057, -12.611684, -0.7244367, 0.18346946, 0.10700805, -107.91296, -13.153835, -0.9124783, 0.12709878, 0.096012175, -101.2308, -13.551485, -1.0773662, 0.07470902, 0.08526665, -94.38393, -13.814306, -1.2199031, 0.026339812, 0.074829005, -87.43731, -13.952125, -1.3409865, -0.018002395, 0.06474949, -80.45097, -13.974832, -1.4415944, -0.058341455, 0.055071317, -73.48, -13.892308, -1.5227703, -0.09472873, 0.04583096, -66.57456, -13.714346, -1.5856107, -0.12724029, 0.03705848, -59.77995, -13.450592, -1.6312516, -0.15597418, 0.028777855, -53.13669, -13.11048, -1.6608567, -0.18104783, 0.021007333},
		'{-1.5015588e-11, 2.1104364e-12, 7.663234e-13, 6.098396e-14, -3.869166e-15, -1.418327e-11, 1.9934542e-12, 7.238459e-13, 5.76036e-14, -3.654697e-15, -1.3397087e-11, 1.8829565e-12, 6.8372294e-13, 5.4410615e-14, -3.452116e-15, -1.26544825e-11, 1.7785837e-12, 6.45824e-13, 5.1394622e-14, -3.2607643e-15, -1.1953041e-11, 1.6799963e-12, 6.1002576e-13, 4.8545803e-14, -3.0800191e-15, -1.1290481e-11, 1.5868736e-12, 5.762119e-13, 4.5854894e-14, -2.9092928e-15, -1.0664646e-11, 1.4989128e-12, 5.442723e-13, 4.3313145e-14, -2.74803e-15, -1.0073502e-11, 1.4158276e-12, 5.1410314e-13, 4.0912284e-14, -2.5957058e-15, -9.515125e-12, 1.3373479e-12, 4.8560624e-13, 3.8644506e-14, -2.4518252e-15, -8.987699e-12, 1.2632184e-12, 4.5868897e-13, 3.650243e-14, -2.3159198e-15, -8.489509e-12, 1.1931978e-12, 4.332637e-13, 3.447909e-14, -2.1875477e-15, -8.018933e-12, 1.1270585e-12, 4.0924778e-13, 3.2567905e-14, -2.0662913e-15, -7.574441e-12, 1.0645854e-12, 3.8656304e-13, 3.0762658e-14, -1.9517562e-15, -7.1545873e-12, 1.0055751e-12, 3.6513576e-13, 2.9057475e-14, -1.8435698e-15, -6.7580065e-12, 9.498358e-13, 3.4489618e-13, 2.744681e-14, -1.7413803e-15, -6.3834086e-12, 8.971861e-13, 3.257785e-13, 2.5925425e-14, -1.6448551e-15, -6.0295744e-12, 8.474548e-13, 3.0772048e-13, 2.4488373e-14, -1.5536802e-15, -5.6953535e-12, 8.004802e-13, 2.9066346e-13, 2.3130976e-14, -1.4675593e-15, -5.379658e-12, 7.561093e-13, 2.745519e-13, 2.1848818e-14, -1.3862121e-15, -5.081462e-12, 7.1419796e-13, 2.593334e-13, 2.0637732e-14, -1.309374e-15, -4.7997955e-12, 6.746098e-13, 2.4495849e-13, 1.9493777e-14, -1.236795e-15, -4.5337414e-12, 6.37216e-13, 2.3138037e-13, 1.841323e-14, -1.1682392e-15, -4.282435e-12, 6.018949e-13, 2.185549e-13, 1.7392582e-14, -1.1034833e-15, -4.045058e-12, 5.685317e-13, 2.0644033e-13, 1.6428506e-14, -1.0423169e-15, -3.8208395e-12, 5.3701786e-13, 1.9499728e-13, 1.5517869e-14, -9.84541e-16}};
	localparam real hf[0:1499] = {0.041534796, -0.00025106283, -0.00029157574, 2.7978147e-06, 5.82289e-06, 0.041284204, -0.00075033685, -0.00028448508, 8.326207e-06, 5.687937e-06, 0.040785868, -0.0012411007, -0.00027042086, 1.3654857e-05, 5.4220955e-06, 0.040045436, -0.0017178204, -0.00024961328, 1.8656523e-05, 5.033122e-06, 0.03907127, -0.0021751644, -0.00022240085, 2.321193e-05, 4.5320057e-06, 0.037874334, -0.0026080792, -0.00018922379, 2.7212154e-05, 3.932477e-06, 0.03646804, -0.0030118593, -0.00015061545, 3.0560703e-05, 3.2505068e-06, 0.034868043, -0.0033822125, -0.000107192514, 3.317523e-05, 2.5037984e-06, 0.033092033, -0.0037153156, -5.9643706e-05, 3.498891e-05, 1.7112812e-06, 0.031159483, -0.004007865, -8.71752e-06, 3.5951427e-05, 8.926147e-07, 0.029091382, -0.004257118, 4.4790846e-05, 3.6029665e-05, 6.7710374e-08, 0.02690994, -0.0044609215, 0.00010005313, 3.520796e-05, -7.4372235e-07, 0.024638291, -0.0046177385, 0.0001562219, 3.348807e-05, -1.5226002e-06, 0.022300186, -0.0047266576, 0.0002124445, 3.08888e-05, -2.2508545e-06, 0.019919666, -0.004787397, 0.00026787687, 2.7445309e-05, -2.9117798e-06, 0.017520765, -0.004800299, 0.00032169677, 2.3208151e-05, -3.4903378e-06, 0.015127185, -0.004766313, 0.00037311652, 1.8242059e-05, -3.9734164e-06, 0.012762014, -0.004686971, 0.00042139483, 1.2624505e-05, -4.3500386e-06, 0.0104474295, -0.0045643575, 0.00046584764, 6.4440724e-06, -4.611522e-06, 0.00820444, -0.0044010663, 0.00050585775, -2.0132107e-07, -4.751589e-06, 0.0060526365, -0.004200157, 0.0005408832, -7.206319e-06, -4.766427e-06, 0.0040099784, -0.0039650984, 0.0005704643, -1.44601e-05, -4.654699e-06, 0.002092596, -0.0036997166, 0.0005942291, -2.1848395e-05, -4.4175094e-06, 0.00031463295, -0.0034081284, 0.00061189727, -2.9255505e-05, -4.058328e-06, -0.0013118859, -0.0030946804, 0.0006232827, -3.6566307e-05, -3.582867e-06, -0.0027771527, -0.0027638816, 0.0006282943, -4.3668166e-05, -2.9989294e-06, -0.004073641, -0.0024203376, 0.0006269355, -5.0452807e-05, -2.3162183e-06, -0.005196136, -0.0020686835, 0.0006193019, -5.6817997e-05, -1.5461219e-06, -0.006141737, -0.0017135186, 0.0006055781, -6.2669154e-05, -7.014739e-07, -0.0069098184, -0.0013593443, 0.00058603287, -6.792074e-05, 2.0370419e-07, -0.007501969, -0.0010105032, 0.000561013, -7.249747e-05, 1.1544739e-06, -0.007921898, -0.0006711236, 0.0005309366, -7.6335375e-05, 2.135259e-06, -0.0081753135, -0.00034506852, 0.00049628475, -7.9382575e-05, 3.130127e-06, -0.008269779, -3.5888985e-05, 0.00045759339, -8.1599894e-05, 4.1230696e-06, -0.008214549, 0.00025321555, 0.0004154435, -8.296122e-05, 5.0982767e-06, -0.00802038, 0.0005194313, 0.00037045157, -8.345366e-05, 6.0403986e-06, -0.0076993345, 0.0007603575, 0.00032325956, -8.3077495e-05, 6.9347943e-06, -0.007264567, 0.0009740267, 0.00027452473, -8.184589e-05, 7.7677605e-06, -0.006730106, 0.0011589184, 0.00022490944, -7.978439e-05, 8.526739e-06, -0.0061106253, 0.0013139657, 0.00017507143, -7.693034e-05, 9.200501e-06, -0.0054212194, 0.001438555, 0.00012565407, -7.3331976e-05, 9.779301e-06, -0.0046771774, 0.0015325192, 7.7277364e-05, -6.9047506e-05, 1.0255004e-05, -0.003893763, 0.0015961247, 3.052947e-05, -6.414397e-05, 1.0621186e-05, -0.003086002, 0.0016300521, -1.4041071e-05, -5.8696005e-05, 1.0873203e-05, -0.0022684818, 0.0016353722, -5.5932254e-05, -5.2784588e-05, 1.1008219e-05, -0.0014551623, 0.0016135158, -9.469464e-05, -4.649562e-05, 1.1025223e-05, -0.00065920514, 0.001566241, -0.00012993641, -3.9918534e-05, 1.0924999e-05, 0.00010718096, 0.0014955952, -0.00016132742, -3.3144854e-05, 1.0710076e-05, 0.0008328751, 0.0014038746, -0.00018860218, -2.6266784e-05, 1.0384654e-05, 0.0015079578, 0.0012935818, -0.00021156181, -1.9375813e-05, 9.954496e-06, 0.0021238036, 0.0011673816, -0.0002300749, -1.2561353e-05, 9.426808e-06, 0.00267315, 0.0010280559, -0.00024407731, -5.9094777e-06, 8.810093e-06, 0.003150146, 0.0008784578, -0.00025357108, 4.9827673e-07, 8.1139915e-06, 0.0035503746, 0.00072146766, -0.0002586222, 6.585999e-06, 7.3491037e-06, 0.0038708579, 0.0005599489, -0.00025935765, 1.2284375e-05, 6.526811e-06, 0.004110036, 0.00039670657, -0.00025596155, 1.753153e-05, 5.659079e-06, 0.0042677284, 0.0002344476, -0.00024867058, 2.2273744e-05, 4.758265e-06, 0.004345076, 7.574436e-05, -0.0002377687, 2.6465998e-05, 3.8369194e-06, 0.0043444666, -7.6998505e-05, -0.00022358146, 3.007241e-05, 2.9075927e-06, 0.0042694397, -0.00022157375, -0.00020646975, 3.306648e-05, 1.9826468e-06, 0.0041245855, -0.00035599695, -0.00018682326, 3.5431218e-05, 1.0740738e-06, 0.003915426, -0.0004785277, -0.00016505376, 3.71591e-05, 1.9332649e-07, 0.0036482878, -0.0005876865, -0.00014158816, 3.8251907e-05, -6.4883864e-07, 0.0033301709, -0.0006822667, -0.00011686175, 3.872039e-05, -1.442503e-06, 0.002968607, -0.0007613425, -9.131136e-05, 3.858387e-05, -2.178711e-06, 0.0025715213, -0.0008242718, -6.53688e-05, 3.7869646e-05, -2.849576e-06, 0.0021470883, -0.00087069476, -3.9454615e-05, 3.661237e-05, -3.4483685e-06, 0.0017035934, -0.00090052845, -1.3972208e-05, 3.4853285e-05, -3.969582e-06, 0.001249296, -0.00091395725, 1.06976095e-05, 3.263941e-05, -4.4089807e-06, 0.0007922993, -0.00091141934, 3.420151e-05, 3.0022655e-05, -4.763623e-06, 0.00034042718, -0.00089359016, 5.621796e-05, 2.705888e-05, -5.0318704e-06, -9.888928e-05, -0.0008613626, 7.646092e-05, 2.3806966e-05, -5.213369e-06, -0.00051871524, -0.0008158246, 9.468285e-05, 2.0327805e-05, -5.3090184e-06, -0.0009127036, -0.00075823476, 0.00011067708, 1.6683356e-05, -5.3209187e-06, -0.0012751736, -0.00068999594, 0.0001242794, 1.2935674e-05, -5.2523037e-06, -0.0016011767, -0.0006126279, 0.000135369, 9.145986e-06, -5.107456e-06, -0.001886547, -0.00052773894, 0.00014386876, 5.3738077e-06, -4.891611e-06, -0.0021279391, -0.00043699733, 0.00014974474, 1.6761131e-06, -4.610849e-06, -0.0023228514, -0.00034210266, 0.00015300514, -1.8934277e-06, -4.2719776e-06, -0.002469633, -0.00024475812, 0.00015369864, -5.285136e-06, -3.8824082e-06, -0.0025674808, -0.0001466433, 0.00015191213, -8.45393e-06, -3.450024e-06, -0.0026164197, -4.9388746e-05, 0.00014776793, -1.1359837e-05, -2.983049e-06, -0.0026172728, 4.544807e-05, 0.0001414207, -1.3968416e-05, -2.4899134e-06, -0.0025716187, 0.00013640465, 0.00013305375, -1.6251079e-05, -1.9791212e-06, -0.00248174, 0.00022213308, 0.00012287522, -1.8185305e-05, -1.4591213e-06, -0.0023505604, 0.00030141728, 0.000111113935, -1.9754776e-05, -9.3818284e-07, -0.0021815759, 0.00037318736, 9.801511e-05, -2.094939e-05, -4.2427752e-07, -0.0019787785, 0.00043653135, 8.383593e-05, -2.176519e-05, 7.502879e-08, -0.0017465743, 0.000490704, 6.884111e-05, -2.220421e-05, 5.526759e-07, -0.0014896997, 0.00053513265, 5.329856e-05, -2.2274216e-05, 1.0021976e-06, -0.0012131332, 0.00056942005, 3.7475045e-05, -2.1988382e-05, 1.4177976e-06, -0.0009220082, 0.0005933447, 2.1632093e-05, -2.1364898e-05, 1.7944142e-06, -0.0006215252, 0.00060685794, 6.0221128e-06, -2.0426502e-05, 2.1277697e-06, -0.00031686708, 0.000610079, -9.115222e-06, -1.9199964e-05, 2.4144072e-06, -1.3116588e-05, 0.0006032868, -2.3556257e-05, -1.771554e-05, 2.6517146e-06, 0.00028482094, 0.0005869106, -3.709627e-05, -1.6006365e-05, 2.8379332e-06, 0.0005722898, 0.0005615176, -4.9552003e-05, -1.4107845e-05, 2.9721539e-06, 0.0008449497, 0.0005277994, -6.076376e-05, -1.2057032e-05, 3.0543008e-06, 0.001098834, 0.000486557, -7.059706e-05, -9.891985e-06, 3.085102e-06, 0.0013304005, 0.00043868393, -7.894386e-05, -7.651149e-06, 3.06605e-06, 0.0015365733, 0.00038514961, -8.572333e-05, -5.3727435e-06, 2.9993512e-06, 0.0017147767, 0.00032698113, -9.088212e-05, -3.094183e-06, 2.8878662e-06, 0.0018629591, 0.00026524524, -9.439426e-05, -8.515203e-07, 2.7350422e-06, 0.001979608, 0.00020103023, -9.626061e-05, 1.3210607e-06, 2.5448396e-06, 0.0020637577, 0.00013542802, -9.650791e-05, 3.3917102e-06, 2.321652e-06, 0.0021149844, 6.951695e-05, -9.518744e-05, 5.331324e-06, 2.070223e-06, 0.0021333976, 4.3451932e-06, -9.237341e-05, 7.113898e-06, 1.795561e-06, 0.0021196199, -5.908462e-05, -8.816096e-05, 8.716823e-06, 1.502852e-06, 0.0020747606, -0.000119829674, -8.266398e-05, 1.0121115e-05, 1.1973733e-06, 0.002000383, -0.00017701974, -7.6012664e-05, 1.1311585e-05, 8.844084e-07, 0.0018984649, -0.00022986843, -6.835092e-05, 1.2276939e-05, 5.691655e-07, 0.0017713541, -0.00027768273, -5.9833645e-05, 1.3009816e-05, 2.5669905e-07, 0.0016217204, -0.00031987083, -5.0623927e-05, 1.35067685e-05, -4.8162583e-08, 0.0014525024, -0.00035594788, -4.089022e-05, 1.3768174e-05, -3.408843e-07, 0.001266854, -0.00038554022, -3.0803512e-05, 1.3798097e-05, -6.1728406e-07, 0.0010680873, -0.00040838748, -2.0534582e-05, 1.3604099e-05, -8.7358524e-07, 0.0008596161, -0.0004243429, -1.0251324e-05, 1.3196993e-05, -1.106461e-06, 0.0006448997, -0.00043337187, -1.1622957e-07, 1.2590566e-05, -1.3130701e-06, 0.00042738713, -0.0004355489, 9.715975e-06, 1.180126e-05, -1.4910838e-06, 0.00021046394, -0.00043105264, 1.9100476e-05, 1.0847818e-05, -1.6387039e-06, -2.5985123e-06, -0.00042015998, 2.7904307e-05, 9.750918e-06, -1.7546723e-06, -0.00020869027, -0.00040323817, 3.600802e-05, 8.532781e-06, -1.8382717e-06, -0.00040490585, -0.00038073648, 4.3307093e-05, 7.216767e-06, -1.8893174e-06, -0.0005885828, -0.00035317618, 4.9713064e-05, 5.8269757e-06, -1.9081417e-06, -0.00075733534, -0.0003211403, 5.515437e-05, 4.387843e-06, -1.8955704e-06, -0.0009090821, -0.00028526245, 5.9576894e-05, 2.923747e-06, -1.8528937e-06, -0.0010420689, -0.00024621532, 6.2944215e-05, 1.4586296e-06, -1.7818282e-06, -0.0011548854, -0.00020469894, 6.523761e-05, 1.5637731e-08, -1.6844771e-06, -0.0012464753, -0.0001614289, 6.645571e-05, -1.3832115e-06, -1.5632824e-06, -0.0013161416, -0.00011712479, 6.661398e-05, -2.7173355e-06, -1.4209761e-06, -0.0013635461, -7.249879e-05, 6.5743894e-05, -3.9678594e-06, -1.2605273e-06, -0.0013887023, -2.8244982e-05, 6.3891915e-05, -5.117852e-06, -1.0850872e-06, -0.001391964, 1.4970881e-05, 6.111827e-05, -6.152525e-06, -8.9793434e-07, -0.0013740092, 5.652074e-05, 5.749555e-05, -7.05939e-06, -7.024187e-07, -0.0013358181, 9.582273e-05, 5.3107167e-05, -7.8283765e-06, -5.0190675e-07, -0.0012786493, 0.00013234868, 4.8045702e-05, -8.451907e-06, -2.997288e-07, -0.0012040103, 0.00016563048, 4.241116e-05, -8.92493e-06, -9.9127995e-08, -0.001113627, 0.00019526538, 3.6309157e-05, -9.2449145e-06, 9.678735e-08, -0.0010094087, 0.0002209201, 2.9849096e-05, -9.411807e-06, 2.850875e-07, -0.0008934142, 0.00024233363, 2.3142342e-05, -9.427944e-06, 4.6306107e-07, -0.0007678137, 0.00025931885, 1.6300424e-05, -9.297936e-06, 6.282498e-07, -0.00063485274, 0.00027176307, 9.433303e-06, -9.028526e-06, 7.7847824e-07, -0.00049681455, 0.0002796273, 2.6477057e-06, -8.628403e-06, 9.118783e-07, -0.0003559839, 0.0002829443, -3.954416e-06, -8.108007e-06, 1.0269079e-06, -0.00021461176, 0.0002818158, -1.0277314e-05, -7.4793093e-06, 1.1223634e-06, -7.4881806e-05, 0.00027640862, -1.6232718e-05, -6.755569e-06, 1.1973882e-06, 6.112102e-05, 0.00026694988, -2.1740963e-05, -5.951088e-06, 1.251473e-06, 0.00019143926, 0.00025372155, -2.6731934e-05, -5.0809535e-06, 1.2844527e-06, 0.00031426887, 0.00023705418, -3.114583e-05, -4.1607746e-06, 1.2964974e-06, 0.00042798184, 0.00021732027, -3.493377e-05, -3.2064231e-06, 1.2880981e-06, 0.0005311455, 0.0001949271, -3.805816e-05, -2.2337795e-06, 1.2600486e-06, 0.00062253774, 0.00017030917, -4.0492905e-05, -1.258483e-06, 1.2134229e-06, 0.00070115924, 0.00014392076, -4.222345e-05, -2.9569895e-07, 1.1495486e-06, 0.0007662408, 0.00011622807, -4.32466e-05, 6.4010254e-07, 1.0699782e-06, 0.00081724813, 8.770176e-05, -4.35702e-05, 1.5353475e-06, 9.764574e-07, 0.0008538814, 5.8809463e-05, -4.3212636e-05, 2.377539e-06, 8.708911e-07, 0.00087607274, 3.0008674e-05, -4.2202217e-05, 3.1554157e-06, 7.553087e-07, 0.00088397873, 1.7400338e-06, -4.0576382e-05, 3.859085e-06, 6.318283e-07, 0.00087797106, -2.5578918e-05, -3.8380836e-05, 4.480132e-06, 5.0262054e-07, 0.000858623, -5.155941e-05, -3.5668552e-05, 5.011698e-06, 3.6987356e-07, 0.000826694, -7.584648e-05, -3.249872e-05, 5.4485395e-06, 2.3575794e-07, 0.0007831117, -9.812332e-05, -2.8935612e-05, 5.7870507e-06, 1.0239382e-07, 0.0007289518, -0.00011811488, -2.504742e-05, 6.0252696e-06, -2.8180478e-08, 0.0006654164, -0.00013559072, -2.0905076e-05, 6.162849e-06, -1.5403734e-07, 0.00059381133, -0.00015036705, -1.6581056e-05, 6.2010117e-06, -2.7338612e-07, 0.00051552226, -0.00016230803, -1.214821e-05, 6.1424766e-06, -3.8459638e-07, 0.00043199077, -0.0001713262, -7.678622e-06, 5.9913687e-06, -4.862178e-07, 0.0003446901, -0.00017738224, -3.2425198e-06, 5.753106e-06, -5.7699685e-07, 0.00025510127, -0.00018048396, 1.0927498e-06, 5.434275e-06, -6.558894e-07, 0.00016469005, -0.00018068451, 5.263664e-06, 5.0424865e-06, -7.220701e-07, 7.488465e-05, -0.0001780801, 9.21138e-06, 4.5862266e-06, -7.74938e-07, -1.2944907e-05, -0.00017280705, 1.2882487e-05, 4.0746936e-06, -8.141181e-07, -9.750609e-05, -0.0001650383, 1.622965e-05, 3.5176333e-06, -8.3945974e-07, -0.00017760119, -0.00015497948, 1.9212137e-05, 2.9251694e-06, -8.510316e-07, -0.0002521426, -0.0001428647, 2.179623e-05, 2.307633e-06, -8.49113e-07, -0.0003201659, -0.00012895184, 2.3955507e-05, 1.6753972e-06, -8.341828e-07, -0.00038084065, -0.00011351787, 2.5671005e-05, 1.0387151e-06, -8.0690523e-07, -0.00043347856, -9.685387e-05, 2.6931266e-05, 4.0756368e-07, -7.6811324e-07, -0.00047753938, -7.926006e-05, 2.7732256e-05, -2.0849993e-07, -7.1879026e-07, -0.00051263423, -6.104082e-05, 2.8077182e-05, -8.004729e-07, -6.600497e-07, -0.00053852645, -4.2499843e-05, 2.7976193e-05, -1.3600273e-06, -5.931133e-07, -0.0005551301, -2.3935505e-05, 2.7445998e-05, -1.8796164e-06, -5.1928896e-07, -0.0005625061, -5.6363674e-06, 2.6509371e-05, -2.3525652e-06, -4.399471e-07, -0.0005608564, 1.2122926e-05, 2.5194613e-05, -2.773144e-06, -3.5649768e-07, -0.000550516, 2.9085437e-05, 2.3534907e-05, -3.136626e-06, -2.7036694e-07, -0.00053194317, 4.5015313e-05, 2.1567657e-05, -3.4393265e-06, -1.829748e-07, -0.0005057082, 5.970072e-05, 1.9333756e-05, -3.6786248e-06, -9.571304e-08, -0.0004724809, 7.29563e-05, 1.6876844e-05, -3.8529683e-06, -9.924751e-09, -0.00043301654, 8.4625186e-05, 1.4242524e-05, -3.961862e-06, 7.311487e-08, -0.00038814152, 9.4580384e-05, 1.1477609e-05, -4.0058394e-06, 1.5221593e-07, -0.000338738, 0.00010272581, 8.629347e-06, -3.98642e-06, 2.2628946e-07, -0.00028572837, 0.0001089967, 5.744669e-06, -3.9060515e-06, 2.943608e-07, -0.00023005955, 0.00011335952, 2.8694867e-06, -3.768044e-06, 3.555809e-07, -0.00017268756, 0.00011581148, 4.8004853e-08, -3.5764851e-06, 4.0923527e-07, -0.0001145623, 0.00011637951, -2.6779e-06, -3.3361537e-06, 4.547504e-07, -5.6613084e-05, 0.00011511882, -5.269251e-06, -3.0524216e-06, 4.9169796e-07, 2.650982e-07, 0.0001121111, -7.690474e-06, -2.7311503e-06, 5.197967e-07, 5.522427e-05, 0.000107462365, -9.90984e-06, -2.3785838e-06, 5.389114e-07, 0.00010747505, 0.00010130049, -1.1899816e-05, -2.0012399e-06, 5.4905075e-07, 0.00015629685, 9.377246e-05, -1.3637359e-05, -1.6057982e-06, 5.503617e-07, 0.00020104682, 8.504147e-05, -1.5104117e-05, -1.1989931e-06, 5.431227e-07, 0.00024116704, 7.5283846e-05, -1.628655e-05, -7.875069e-07, 5.277355e-07, 0.00027619046, 6.4685846e-05, -1.7175993e-05, -3.7786796e-07, 5.0471385e-07, 0.00030574488, 5.344045e-05, -1.7768598e-05, 2.3644843e-08, 4.746725e-07, 0.00032955565, 4.1744155e-05, -1.806526e-05, 4.11091e-07, 4.3831406e-07, 0.0003474466, 2.9793786e-05, -1.8071425e-05, 7.7894896e-07, 3.964151e-07, 0.00035933938, 1.7783444e-05, -1.7796852e-05, 1.1221874e-06, 3.4981156e-07, 0.0003652514, 5.9015915e-06, -1.7255326e-05, 1.4363266e-06, 2.993841e-07, 0.0003652924, -5.671682e-06, -1.6464299e-05, 1.717489e-06, 2.460427e-07, 0.0003596594, -1.6767168e-05, -1.5444495e-05, 1.9624395e-06, 1.9071163e-07, 0.0003486309, -2.7228793e-05, -1.42194895e-05, 2.1686124e-06, 1.3431476e-07, 0.0003325598, -3.6915593e-05, -1.2815233e-05, 2.3341308e-06, 7.776114e-08, 0.00031186524, -4.5703397e-05, -1.1259582e-05, 2.4578098e-06, 2.1931545e-08, 0.000287024, -5.3486165e-05, -9.5817895e-06, 2.5391537e-06, -3.23343e-08, 0.00025856117, -6.017704e-05, -7.812017e-06, 2.5783388e-06, -8.424928e-08, 0.00022704026, -6.570903e-05, -5.9808294e-06, 2.5761885e-06, -1.3308932e-07, 0.00019305323, -7.003539e-05, -4.1187063e-06, 2.5341392e-06, -1.7820247e-07, 0.00015721038, -7.3129646e-05, -2.255579e-06, 2.454196e-06, -2.1901654e-07, 0.00012013018, -7.498532e-05, -4.2037928e-07, 2.3388839e-06, -2.550453e-07, 8.242948e-05, -7.56154e-05, 1.3593717e-06, 2.19119e-06, -2.858931e-07, 4.4713957e-05, -7.505139e-05, 3.057944e-06, 2.0145026e-06, -3.1125788e-07, 7.5691023e-06, -7.3342286e-05, 4.6517366e-06, 1.8125437e-06, -3.3093275e-07, -2.8448172e-05, -7.0553186e-05, 6.1195706e-06, 1.5893014e-06, -3.4480598e-07, -6.2817206e-05, -6.676372e-05, 7.4429367e-06, 1.3489584e-06, -3.5285944e-07, -9.506044e-05, -6.206637e-05, 8.606192e-06, 1.0958212e-06, -3.5516578e-07, -0.00012474938, -5.6564564e-05, 9.596702e-06, 8.342483e-07, -3.5188424e-07, -0.00015150955, -5.037071e-05, 1.040494e-05, 5.6858164e-07, -3.4325524e-07, -0.00017502453, -4.3604156e-05, 1.1024528e-05, 3.0307976e-07, -3.2959383e-07, -0.00019503887, -3.6389116e-05, 1.1452226e-05, 4.185431e-08, -3.112825e-07, -0.00021135999, -2.8852557e-05, 1.168788e-05, -2.1118834e-07, -2.8876266e-07, -0.00022385905, -2.1122156e-05, 1.1734318e-05, -4.5240088e-07, -2.6252616e-07, -0.00023247086, -1.3324285e-05, 1.1597205e-05, -6.7844275e-07, -2.3310567e-07, -0.0002371926, -5.5821024e-06, 1.1284865e-05, -8.8632163e-07, -2.0106522e-07, -0.00023808192, 1.9862475e-06, 1.080805e-05, -1.0734279e-06, -1.6699035e-07, -0.00023525392, 9.269301e-06, 1.0179707e-05, -1.2375623e-06, -1.3147829e-07, -0.00022887741, 1.6163774e-05, 9.414689e-06, -1.3769558e-06, -9.512833e-08, -0.00021917057, 2.257589e-05, 8.529469e-06, -1.4902831e-06, -5.8532482e-08, -0.00020639582, 2.842251e-05, 7.541826e-06, -1.5766676e-06, -2.226652e-08, -0.0001908543, 3.3632063e-05, 6.4705287e-06, -1.6356801e-06, 1.311837e-08, -0.0001728799, 3.8145266e-05, 5.335007e-06, -1.6673299e-06, 4.7103306e-08, -0.00015283293, 4.191563e-05, 4.155031e-06, -1.6720508e-06, 7.920866e-08, -0.00013109372, 4.4909746e-05, 2.950394e-06, -1.6506789e-06, 1.0900016e-07, -0.00010805603, 4.7107358e-05, 1.7406019e-06, -1.6044269e-06, 1.360941e-07, -8.4120424e-05, 4.8501246e-05, 5.4458303e-07, -1.5348518e-06, 1.6016155e-07, -5.968793e-05, 4.9096885e-05, -6.195867e-07, -1.4438201e-06, 1.8093162e-07, -3.5153746e-05, 4.8911937e-05, -1.734935e-06, -1.3334676e-06, 1.9819372e-07, -1.09013345e-05, 4.797557e-05, -2.7858193e-06, -1.2061573e-06, 2.117987e-07, 1.27031235e-05, 4.6327605e-05, -3.7581237e-06, -1.0644358e-06, 2.2165922e-07, 3.531583e-05, 4.401756e-05, -4.639427e-06, -9.109866e-07, 2.2774888e-07, 5.6619927e-05, 4.1103536e-05, -5.4191373e-06, -7.485846e-07, 2.3010065e-07, 7.632953e-05, 3.7651036e-05, -6.088595e-06, -5.8004986e-07, 2.2880432e-07, 9.419308e-05, 3.37317e-05, -6.6411417e-06, -4.082021e-07, 2.2400322e-07, 0.0001099961, 2.9421984e-05, -7.0721553e-06, -2.3581738e-07, 2.1589014e-07, 0.00012356327, 2.4801822e-05, -7.379054e-06, -6.5586256e-08, 2.0470272e-07, 0.0001347598, 1.9953257e-05, -7.5612647e-06, 9.992489e-08, 1.9071823e-07, 0.00014349222, 1.4959106e-05, -7.6201695e-06, 2.5830948e-07, 1.7424792e-07, 0.00014970833, 9.901651e-06, -7.5590124e-06, 4.0735262e-07, 1.5563107e-07, 0.00015339672, 4.861377e-06, -7.3827896e-06, 5.45059e-07, 1.3522879e-07, 0.00015458548, -8.420873e-08, -7.098112e-06, 6.6967635e-07, 1.1341764e-07, 0.00015334053, -4.861681e-06, -6.7130477e-06, 7.7971447e-07, 9.058333e-08, 0.00014976322, -9.402696e-06, -6.23695e-06, 8.739594e-07, 6.711439e-08, 0.00014398767, -1.364488e-05, -5.680266e-06, 9.514829e-07, 4.339609e-08, 0.00013617745, -1.7532591e-05, -5.05434e-06, 1.0116473e-06, 1.9804533e-08, 0.00012652224, -2.1017559e-05, -4.371206e-06, 1.0541056e-06, -3.2988252e-09, 0.0001152338, -2.4059378e-05, -3.6433796e-06, 1.0787968e-06, -2.5572303e-08, 0.00010254213, -2.662588e-05, -2.8836455e-06, 1.0859374e-06, -4.669862e-08, 8.869116e-05, -2.8693334e-05, -2.1048527e-06, 1.0760084e-06, -6.638898e-08, 7.393456e-05, -3.0246556e-05, -1.3197115e-06, 1.0497396e-06, -8.43866e-08, 5.853149e-05, -3.127883e-05, -5.406018e-07, 1.008089e-06, -1.0046959e-07, 4.274236e-05, -3.1791744e-05, 2.2060745e-07, 9.522209e-07, -1.1445326e-07, 2.6824775e-05, -3.1794883e-05, 9.527252e-07, 8.834806e-07, -1.2619164e-07, 1.1029648e-05, -3.1305397e-05, 1.6453887e-06, 8.0336747e-07, -1.3557855e-07, -4.402484e-06, -3.0347495e-05, 2.2891963e-06, 7.1350655e-07, -1.4254776e-07, -1.9244822e-05, -2.8951832e-05, 2.8758209e-06, 6.156193e-07, -1.4707284e-07, -3.328736e-05, -2.7154802e-05, 3.3981019e-06, 5.114932e-07, -1.4916608e-07, -4.633957e-05, -2.4997797e-05, 3.8501175e-06, 4.0295237e-07, -1.4887705e-07, -5.8232705e-05, -2.2526383e-05, 4.2272345e-06, 2.9182763e-07, -1.4629057e-07, -6.882166e-05, -1.9789464e-05, 4.5261377e-06, 1.7992816e-07, -1.4152423e-07, -7.7986435e-05, -1.6838409e-05, 4.7448334e-06, 6.901412e-08, -1.3472541e-07, -8.563317e-05, -1.3726165e-05, 4.8826405e-06, -3.922905e-08, -1.2606803e-07, -9.169465e-05, -1.0506393e-05, 4.9401533e-06, -1.4321412e-07, -1.15748946e-07, -9.613054e-05, -7.2326084e-06, 4.919189e-06, -2.4147343e-07, -1.0398412e-07, -9.8927005e-05, -3.9573574e-06, 4.8227216e-06, -3.3267753e-07, -9.100465e-08, -0.00010009611, -7.314347e-07, 4.654794e-06, -4.156512e-07, -7.705263e-08, -9.967471e-05, 2.3968441e-06, 4.4204185e-06, -4.8938637e-07, -6.237709e-08, -9.7723074e-05, 5.382307e-06, 4.12547e-06, -5.5305213e-07, -4.722985e-08, -9.432313e-05, 8.18352e-06, 3.7765624e-06, -6.060018e-07, -3.1861553e-08, -8.957648e-05, 1.0763302e-05, 3.3809233e-06, -6.4777635e-07, -1.6517804e-08, -8.360217e-05, 1.3089159e-05, 2.9462597e-06, -6.7810555e-07, -1.4355486e-09, -7.653425e-05, 1.5133629e-05, 2.4806236e-06, -6.969056e-07, 1.316032e-08, -6.851917e-05, 1.6874536e-05, 1.9922754e-06, -7.0427427e-07, 2.7060032e-08, -5.9713133e-05, 1.8295155e-05, 1.489548e-06, -7.00483e-07, 4.0071686e-08, -5.0279305e-05, 1.9384292e-05, 9.807164e-07, -6.859671e-07, 5.2023616e-08, -4.0385075e-05, 2.0136264e-05, 4.738707e-07, -6.6131344e-07, 6.276637e-08, -3.0199322e-05, 2.0550806e-05, -2.320288e-08, -6.2724604e-07, 7.2174274e-08, -1.9889725e-05, 2.063289e-05, -5.031323e-07, -5.8461046e-07, 8.0146584e-08, -9.6202275e-06, 2.039247e-05, -9.5906e-07, -5.343565e-07, 8.66082e-08, 4.5138748e-07, 1.9844165e-05, -1.384732e-06, -4.7751985e-07, 9.1509975e-08, 1.01757305e-05, 1.900687e-05, -1.7745737e-06, -4.1520332e-07, 9.482858e-08, 1.941384e-05, 1.7903314e-05, -2.1237545e-06, -3.4855745e-07, 9.6566005e-08};
	localparam real hb[0:1499] = {0.041534796, 0.00025106283, -0.00029157574, -2.7978147e-06, 5.82289e-06, 0.041284204, 0.00075033685, -0.00028448508, -8.326207e-06, 5.687937e-06, 0.040785868, 0.0012411007, -0.00027042086, -1.3654857e-05, 5.4220955e-06, 0.040045436, 0.0017178204, -0.00024961328, -1.8656523e-05, 5.033122e-06, 0.03907127, 0.0021751644, -0.00022240085, -2.321193e-05, 4.5320057e-06, 0.037874334, 0.0026080792, -0.00018922379, -2.7212154e-05, 3.932477e-06, 0.03646804, 0.0030118593, -0.00015061545, -3.0560703e-05, 3.2505068e-06, 0.034868043, 0.0033822125, -0.000107192514, -3.317523e-05, 2.5037984e-06, 0.033092033, 0.0037153156, -5.9643706e-05, -3.498891e-05, 1.7112812e-06, 0.031159483, 0.004007865, -8.71752e-06, -3.5951427e-05, 8.926147e-07, 0.029091382, 0.004257118, 4.4790846e-05, -3.6029665e-05, 6.7710374e-08, 0.02690994, 0.0044609215, 0.00010005313, -3.520796e-05, -7.4372235e-07, 0.024638291, 0.0046177385, 0.0001562219, -3.348807e-05, -1.5226002e-06, 0.022300186, 0.0047266576, 0.0002124445, -3.08888e-05, -2.2508545e-06, 0.019919666, 0.004787397, 0.00026787687, -2.7445309e-05, -2.9117798e-06, 0.017520765, 0.004800299, 0.00032169677, -2.3208151e-05, -3.4903378e-06, 0.015127185, 0.004766313, 0.00037311652, -1.8242059e-05, -3.9734164e-06, 0.012762014, 0.004686971, 0.00042139483, -1.2624505e-05, -4.3500386e-06, 0.0104474295, 0.0045643575, 0.00046584764, -6.4440724e-06, -4.611522e-06, 0.00820444, 0.0044010663, 0.00050585775, 2.0132107e-07, -4.751589e-06, 0.0060526365, 0.004200157, 0.0005408832, 7.206319e-06, -4.766427e-06, 0.0040099784, 0.0039650984, 0.0005704643, 1.44601e-05, -4.654699e-06, 0.002092596, 0.0036997166, 0.0005942291, 2.1848395e-05, -4.4175094e-06, 0.00031463295, 0.0034081284, 0.00061189727, 2.9255505e-05, -4.058328e-06, -0.0013118859, 0.0030946804, 0.0006232827, 3.6566307e-05, -3.582867e-06, -0.0027771527, 0.0027638816, 0.0006282943, 4.3668166e-05, -2.9989294e-06, -0.004073641, 0.0024203376, 0.0006269355, 5.0452807e-05, -2.3162183e-06, -0.005196136, 0.0020686835, 0.0006193019, 5.6817997e-05, -1.5461219e-06, -0.006141737, 0.0017135186, 0.0006055781, 6.2669154e-05, -7.014739e-07, -0.0069098184, 0.0013593443, 0.00058603287, 6.792074e-05, 2.0370419e-07, -0.007501969, 0.0010105032, 0.000561013, 7.249747e-05, 1.1544739e-06, -0.007921898, 0.0006711236, 0.0005309366, 7.6335375e-05, 2.135259e-06, -0.0081753135, 0.00034506852, 0.00049628475, 7.9382575e-05, 3.130127e-06, -0.008269779, 3.5888985e-05, 0.00045759339, 8.1599894e-05, 4.1230696e-06, -0.008214549, -0.00025321555, 0.0004154435, 8.296122e-05, 5.0982767e-06, -0.00802038, -0.0005194313, 0.00037045157, 8.345366e-05, 6.0403986e-06, -0.0076993345, -0.0007603575, 0.00032325956, 8.3077495e-05, 6.9347943e-06, -0.007264567, -0.0009740267, 0.00027452473, 8.184589e-05, 7.7677605e-06, -0.006730106, -0.0011589184, 0.00022490944, 7.978439e-05, 8.526739e-06, -0.0061106253, -0.0013139657, 0.00017507143, 7.693034e-05, 9.200501e-06, -0.0054212194, -0.001438555, 0.00012565407, 7.3331976e-05, 9.779301e-06, -0.0046771774, -0.0015325192, 7.7277364e-05, 6.9047506e-05, 1.0255004e-05, -0.003893763, -0.0015961247, 3.052947e-05, 6.414397e-05, 1.0621186e-05, -0.003086002, -0.0016300521, -1.4041071e-05, 5.8696005e-05, 1.0873203e-05, -0.0022684818, -0.0016353722, -5.5932254e-05, 5.2784588e-05, 1.1008219e-05, -0.0014551623, -0.0016135158, -9.469464e-05, 4.649562e-05, 1.1025223e-05, -0.00065920514, -0.001566241, -0.00012993641, 3.9918534e-05, 1.0924999e-05, 0.00010718096, -0.0014955952, -0.00016132742, 3.3144854e-05, 1.0710076e-05, 0.0008328751, -0.0014038746, -0.00018860218, 2.6266784e-05, 1.0384654e-05, 0.0015079578, -0.0012935818, -0.00021156181, 1.9375813e-05, 9.954496e-06, 0.0021238036, -0.0011673816, -0.0002300749, 1.2561353e-05, 9.426808e-06, 0.00267315, -0.0010280559, -0.00024407731, 5.9094777e-06, 8.810093e-06, 0.003150146, -0.0008784578, -0.00025357108, -4.9827673e-07, 8.1139915e-06, 0.0035503746, -0.00072146766, -0.0002586222, -6.585999e-06, 7.3491037e-06, 0.0038708579, -0.0005599489, -0.00025935765, -1.2284375e-05, 6.526811e-06, 0.004110036, -0.00039670657, -0.00025596155, -1.753153e-05, 5.659079e-06, 0.0042677284, -0.0002344476, -0.00024867058, -2.2273744e-05, 4.758265e-06, 0.004345076, -7.574436e-05, -0.0002377687, -2.6465998e-05, 3.8369194e-06, 0.0043444666, 7.6998505e-05, -0.00022358146, -3.007241e-05, 2.9075927e-06, 0.0042694397, 0.00022157375, -0.00020646975, -3.306648e-05, 1.9826468e-06, 0.0041245855, 0.00035599695, -0.00018682326, -3.5431218e-05, 1.0740738e-06, 0.003915426, 0.0004785277, -0.00016505376, -3.71591e-05, 1.9332649e-07, 0.0036482878, 0.0005876865, -0.00014158816, -3.8251907e-05, -6.4883864e-07, 0.0033301709, 0.0006822667, -0.00011686175, -3.872039e-05, -1.442503e-06, 0.002968607, 0.0007613425, -9.131136e-05, -3.858387e-05, -2.178711e-06, 0.0025715213, 0.0008242718, -6.53688e-05, -3.7869646e-05, -2.849576e-06, 0.0021470883, 0.00087069476, -3.9454615e-05, -3.661237e-05, -3.4483685e-06, 0.0017035934, 0.00090052845, -1.3972208e-05, -3.4853285e-05, -3.969582e-06, 0.001249296, 0.00091395725, 1.06976095e-05, -3.263941e-05, -4.4089807e-06, 0.0007922993, 0.00091141934, 3.420151e-05, -3.0022655e-05, -4.763623e-06, 0.00034042718, 0.00089359016, 5.621796e-05, -2.705888e-05, -5.0318704e-06, -9.888928e-05, 0.0008613626, 7.646092e-05, -2.3806966e-05, -5.213369e-06, -0.00051871524, 0.0008158246, 9.468285e-05, -2.0327805e-05, -5.3090184e-06, -0.0009127036, 0.00075823476, 0.00011067708, -1.6683356e-05, -5.3209187e-06, -0.0012751736, 0.00068999594, 0.0001242794, -1.2935674e-05, -5.2523037e-06, -0.0016011767, 0.0006126279, 0.000135369, -9.145986e-06, -5.107456e-06, -0.001886547, 0.00052773894, 0.00014386876, -5.3738077e-06, -4.891611e-06, -0.0021279391, 0.00043699733, 0.00014974474, -1.6761131e-06, -4.610849e-06, -0.0023228514, 0.00034210266, 0.00015300514, 1.8934277e-06, -4.2719776e-06, -0.002469633, 0.00024475812, 0.00015369864, 5.285136e-06, -3.8824082e-06, -0.0025674808, 0.0001466433, 0.00015191213, 8.45393e-06, -3.450024e-06, -0.0026164197, 4.9388746e-05, 0.00014776793, 1.1359837e-05, -2.983049e-06, -0.0026172728, -4.544807e-05, 0.0001414207, 1.3968416e-05, -2.4899134e-06, -0.0025716187, -0.00013640465, 0.00013305375, 1.6251079e-05, -1.9791212e-06, -0.00248174, -0.00022213308, 0.00012287522, 1.8185305e-05, -1.4591213e-06, -0.0023505604, -0.00030141728, 0.000111113935, 1.9754776e-05, -9.3818284e-07, -0.0021815759, -0.00037318736, 9.801511e-05, 2.094939e-05, -4.2427752e-07, -0.0019787785, -0.00043653135, 8.383593e-05, 2.176519e-05, 7.502879e-08, -0.0017465743, -0.000490704, 6.884111e-05, 2.220421e-05, 5.526759e-07, -0.0014896997, -0.00053513265, 5.329856e-05, 2.2274216e-05, 1.0021976e-06, -0.0012131332, -0.00056942005, 3.7475045e-05, 2.1988382e-05, 1.4177976e-06, -0.0009220082, -0.0005933447, 2.1632093e-05, 2.1364898e-05, 1.7944142e-06, -0.0006215252, -0.00060685794, 6.0221128e-06, 2.0426502e-05, 2.1277697e-06, -0.00031686708, -0.000610079, -9.115222e-06, 1.9199964e-05, 2.4144072e-06, -1.3116588e-05, -0.0006032868, -2.3556257e-05, 1.771554e-05, 2.6517146e-06, 0.00028482094, -0.0005869106, -3.709627e-05, 1.6006365e-05, 2.8379332e-06, 0.0005722898, -0.0005615176, -4.9552003e-05, 1.4107845e-05, 2.9721539e-06, 0.0008449497, -0.0005277994, -6.076376e-05, 1.2057032e-05, 3.0543008e-06, 0.001098834, -0.000486557, -7.059706e-05, 9.891985e-06, 3.085102e-06, 0.0013304005, -0.00043868393, -7.894386e-05, 7.651149e-06, 3.06605e-06, 0.0015365733, -0.00038514961, -8.572333e-05, 5.3727435e-06, 2.9993512e-06, 0.0017147767, -0.00032698113, -9.088212e-05, 3.094183e-06, 2.8878662e-06, 0.0018629591, -0.00026524524, -9.439426e-05, 8.515203e-07, 2.7350422e-06, 0.001979608, -0.00020103023, -9.626061e-05, -1.3210607e-06, 2.5448396e-06, 0.0020637577, -0.00013542802, -9.650791e-05, -3.3917102e-06, 2.321652e-06, 0.0021149844, -6.951695e-05, -9.518744e-05, -5.331324e-06, 2.070223e-06, 0.0021333976, -4.3451932e-06, -9.237341e-05, -7.113898e-06, 1.795561e-06, 0.0021196199, 5.908462e-05, -8.816096e-05, -8.716823e-06, 1.502852e-06, 0.0020747606, 0.000119829674, -8.266398e-05, -1.0121115e-05, 1.1973733e-06, 0.002000383, 0.00017701974, -7.6012664e-05, -1.1311585e-05, 8.844084e-07, 0.0018984649, 0.00022986843, -6.835092e-05, -1.2276939e-05, 5.691655e-07, 0.0017713541, 0.00027768273, -5.9833645e-05, -1.3009816e-05, 2.5669905e-07, 0.0016217204, 0.00031987083, -5.0623927e-05, -1.35067685e-05, -4.8162583e-08, 0.0014525024, 0.00035594788, -4.089022e-05, -1.3768174e-05, -3.408843e-07, 0.001266854, 0.00038554022, -3.0803512e-05, -1.3798097e-05, -6.1728406e-07, 0.0010680873, 0.00040838748, -2.0534582e-05, -1.3604099e-05, -8.7358524e-07, 0.0008596161, 0.0004243429, -1.0251324e-05, -1.3196993e-05, -1.106461e-06, 0.0006448997, 0.00043337187, -1.1622957e-07, -1.2590566e-05, -1.3130701e-06, 0.00042738713, 0.0004355489, 9.715975e-06, -1.180126e-05, -1.4910838e-06, 0.00021046394, 0.00043105264, 1.9100476e-05, -1.0847818e-05, -1.6387039e-06, -2.5985123e-06, 0.00042015998, 2.7904307e-05, -9.750918e-06, -1.7546723e-06, -0.00020869027, 0.00040323817, 3.600802e-05, -8.532781e-06, -1.8382717e-06, -0.00040490585, 0.00038073648, 4.3307093e-05, -7.216767e-06, -1.8893174e-06, -0.0005885828, 0.00035317618, 4.9713064e-05, -5.8269757e-06, -1.9081417e-06, -0.00075733534, 0.0003211403, 5.515437e-05, -4.387843e-06, -1.8955704e-06, -0.0009090821, 0.00028526245, 5.9576894e-05, -2.923747e-06, -1.8528937e-06, -0.0010420689, 0.00024621532, 6.2944215e-05, -1.4586296e-06, -1.7818282e-06, -0.0011548854, 0.00020469894, 6.523761e-05, -1.5637731e-08, -1.6844771e-06, -0.0012464753, 0.0001614289, 6.645571e-05, 1.3832115e-06, -1.5632824e-06, -0.0013161416, 0.00011712479, 6.661398e-05, 2.7173355e-06, -1.4209761e-06, -0.0013635461, 7.249879e-05, 6.5743894e-05, 3.9678594e-06, -1.2605273e-06, -0.0013887023, 2.8244982e-05, 6.3891915e-05, 5.117852e-06, -1.0850872e-06, -0.001391964, -1.4970881e-05, 6.111827e-05, 6.152525e-06, -8.9793434e-07, -0.0013740092, -5.652074e-05, 5.749555e-05, 7.05939e-06, -7.024187e-07, -0.0013358181, -9.582273e-05, 5.3107167e-05, 7.8283765e-06, -5.0190675e-07, -0.0012786493, -0.00013234868, 4.8045702e-05, 8.451907e-06, -2.997288e-07, -0.0012040103, -0.00016563048, 4.241116e-05, 8.92493e-06, -9.9127995e-08, -0.001113627, -0.00019526538, 3.6309157e-05, 9.2449145e-06, 9.678735e-08, -0.0010094087, -0.0002209201, 2.9849096e-05, 9.411807e-06, 2.850875e-07, -0.0008934142, -0.00024233363, 2.3142342e-05, 9.427944e-06, 4.6306107e-07, -0.0007678137, -0.00025931885, 1.6300424e-05, 9.297936e-06, 6.282498e-07, -0.00063485274, -0.00027176307, 9.433303e-06, 9.028526e-06, 7.7847824e-07, -0.00049681455, -0.0002796273, 2.6477057e-06, 8.628403e-06, 9.118783e-07, -0.0003559839, -0.0002829443, -3.954416e-06, 8.108007e-06, 1.0269079e-06, -0.00021461176, -0.0002818158, -1.0277314e-05, 7.4793093e-06, 1.1223634e-06, -7.4881806e-05, -0.00027640862, -1.6232718e-05, 6.755569e-06, 1.1973882e-06, 6.112102e-05, -0.00026694988, -2.1740963e-05, 5.951088e-06, 1.251473e-06, 0.00019143926, -0.00025372155, -2.6731934e-05, 5.0809535e-06, 1.2844527e-06, 0.00031426887, -0.00023705418, -3.114583e-05, 4.1607746e-06, 1.2964974e-06, 0.00042798184, -0.00021732027, -3.493377e-05, 3.2064231e-06, 1.2880981e-06, 0.0005311455, -0.0001949271, -3.805816e-05, 2.2337795e-06, 1.2600486e-06, 0.00062253774, -0.00017030917, -4.0492905e-05, 1.258483e-06, 1.2134229e-06, 0.00070115924, -0.00014392076, -4.222345e-05, 2.9569895e-07, 1.1495486e-06, 0.0007662408, -0.00011622807, -4.32466e-05, -6.4010254e-07, 1.0699782e-06, 0.00081724813, -8.770176e-05, -4.35702e-05, -1.5353475e-06, 9.764574e-07, 0.0008538814, -5.8809463e-05, -4.3212636e-05, -2.377539e-06, 8.708911e-07, 0.00087607274, -3.0008674e-05, -4.2202217e-05, -3.1554157e-06, 7.553087e-07, 0.00088397873, -1.7400338e-06, -4.0576382e-05, -3.859085e-06, 6.318283e-07, 0.00087797106, 2.5578918e-05, -3.8380836e-05, -4.480132e-06, 5.0262054e-07, 0.000858623, 5.155941e-05, -3.5668552e-05, -5.011698e-06, 3.6987356e-07, 0.000826694, 7.584648e-05, -3.249872e-05, -5.4485395e-06, 2.3575794e-07, 0.0007831117, 9.812332e-05, -2.8935612e-05, -5.7870507e-06, 1.0239382e-07, 0.0007289518, 0.00011811488, -2.504742e-05, -6.0252696e-06, -2.8180478e-08, 0.0006654164, 0.00013559072, -2.0905076e-05, -6.162849e-06, -1.5403734e-07, 0.00059381133, 0.00015036705, -1.6581056e-05, -6.2010117e-06, -2.7338612e-07, 0.00051552226, 0.00016230803, -1.214821e-05, -6.1424766e-06, -3.8459638e-07, 0.00043199077, 0.0001713262, -7.678622e-06, -5.9913687e-06, -4.862178e-07, 0.0003446901, 0.00017738224, -3.2425198e-06, -5.753106e-06, -5.7699685e-07, 0.00025510127, 0.00018048396, 1.0927498e-06, -5.434275e-06, -6.558894e-07, 0.00016469005, 0.00018068451, 5.263664e-06, -5.0424865e-06, -7.220701e-07, 7.488465e-05, 0.0001780801, 9.21138e-06, -4.5862266e-06, -7.74938e-07, -1.2944907e-05, 0.00017280705, 1.2882487e-05, -4.0746936e-06, -8.141181e-07, -9.750609e-05, 0.0001650383, 1.622965e-05, -3.5176333e-06, -8.3945974e-07, -0.00017760119, 0.00015497948, 1.9212137e-05, -2.9251694e-06, -8.510316e-07, -0.0002521426, 0.0001428647, 2.179623e-05, -2.307633e-06, -8.49113e-07, -0.0003201659, 0.00012895184, 2.3955507e-05, -1.6753972e-06, -8.341828e-07, -0.00038084065, 0.00011351787, 2.5671005e-05, -1.0387151e-06, -8.0690523e-07, -0.00043347856, 9.685387e-05, 2.6931266e-05, -4.0756368e-07, -7.6811324e-07, -0.00047753938, 7.926006e-05, 2.7732256e-05, 2.0849993e-07, -7.1879026e-07, -0.00051263423, 6.104082e-05, 2.8077182e-05, 8.004729e-07, -6.600497e-07, -0.00053852645, 4.2499843e-05, 2.7976193e-05, 1.3600273e-06, -5.931133e-07, -0.0005551301, 2.3935505e-05, 2.7445998e-05, 1.8796164e-06, -5.1928896e-07, -0.0005625061, 5.6363674e-06, 2.6509371e-05, 2.3525652e-06, -4.399471e-07, -0.0005608564, -1.2122926e-05, 2.5194613e-05, 2.773144e-06, -3.5649768e-07, -0.000550516, -2.9085437e-05, 2.3534907e-05, 3.136626e-06, -2.7036694e-07, -0.00053194317, -4.5015313e-05, 2.1567657e-05, 3.4393265e-06, -1.829748e-07, -0.0005057082, -5.970072e-05, 1.9333756e-05, 3.6786248e-06, -9.571304e-08, -0.0004724809, -7.29563e-05, 1.6876844e-05, 3.8529683e-06, -9.924751e-09, -0.00043301654, -8.4625186e-05, 1.4242524e-05, 3.961862e-06, 7.311487e-08, -0.00038814152, -9.4580384e-05, 1.1477609e-05, 4.0058394e-06, 1.5221593e-07, -0.000338738, -0.00010272581, 8.629347e-06, 3.98642e-06, 2.2628946e-07, -0.00028572837, -0.0001089967, 5.744669e-06, 3.9060515e-06, 2.943608e-07, -0.00023005955, -0.00011335952, 2.8694867e-06, 3.768044e-06, 3.555809e-07, -0.00017268756, -0.00011581148, 4.8004853e-08, 3.5764851e-06, 4.0923527e-07, -0.0001145623, -0.00011637951, -2.6779e-06, 3.3361537e-06, 4.547504e-07, -5.6613084e-05, -0.00011511882, -5.269251e-06, 3.0524216e-06, 4.9169796e-07, 2.650982e-07, -0.0001121111, -7.690474e-06, 2.7311503e-06, 5.197967e-07, 5.522427e-05, -0.000107462365, -9.90984e-06, 2.3785838e-06, 5.389114e-07, 0.00010747505, -0.00010130049, -1.1899816e-05, 2.0012399e-06, 5.4905075e-07, 0.00015629685, -9.377246e-05, -1.3637359e-05, 1.6057982e-06, 5.503617e-07, 0.00020104682, -8.504147e-05, -1.5104117e-05, 1.1989931e-06, 5.431227e-07, 0.00024116704, -7.5283846e-05, -1.628655e-05, 7.875069e-07, 5.277355e-07, 0.00027619046, -6.4685846e-05, -1.7175993e-05, 3.7786796e-07, 5.0471385e-07, 0.00030574488, -5.344045e-05, -1.7768598e-05, -2.3644843e-08, 4.746725e-07, 0.00032955565, -4.1744155e-05, -1.806526e-05, -4.11091e-07, 4.3831406e-07, 0.0003474466, -2.9793786e-05, -1.8071425e-05, -7.7894896e-07, 3.964151e-07, 0.00035933938, -1.7783444e-05, -1.7796852e-05, -1.1221874e-06, 3.4981156e-07, 0.0003652514, -5.9015915e-06, -1.7255326e-05, -1.4363266e-06, 2.993841e-07, 0.0003652924, 5.671682e-06, -1.6464299e-05, -1.717489e-06, 2.460427e-07, 0.0003596594, 1.6767168e-05, -1.5444495e-05, -1.9624395e-06, 1.9071163e-07, 0.0003486309, 2.7228793e-05, -1.42194895e-05, -2.1686124e-06, 1.3431476e-07, 0.0003325598, 3.6915593e-05, -1.2815233e-05, -2.3341308e-06, 7.776114e-08, 0.00031186524, 4.5703397e-05, -1.1259582e-05, -2.4578098e-06, 2.1931545e-08, 0.000287024, 5.3486165e-05, -9.5817895e-06, -2.5391537e-06, -3.23343e-08, 0.00025856117, 6.017704e-05, -7.812017e-06, -2.5783388e-06, -8.424928e-08, 0.00022704026, 6.570903e-05, -5.9808294e-06, -2.5761885e-06, -1.3308932e-07, 0.00019305323, 7.003539e-05, -4.1187063e-06, -2.5341392e-06, -1.7820247e-07, 0.00015721038, 7.3129646e-05, -2.255579e-06, -2.454196e-06, -2.1901654e-07, 0.00012013018, 7.498532e-05, -4.2037928e-07, -2.3388839e-06, -2.550453e-07, 8.242948e-05, 7.56154e-05, 1.3593717e-06, -2.19119e-06, -2.858931e-07, 4.4713957e-05, 7.505139e-05, 3.057944e-06, -2.0145026e-06, -3.1125788e-07, 7.5691023e-06, 7.3342286e-05, 4.6517366e-06, -1.8125437e-06, -3.3093275e-07, -2.8448172e-05, 7.0553186e-05, 6.1195706e-06, -1.5893014e-06, -3.4480598e-07, -6.2817206e-05, 6.676372e-05, 7.4429367e-06, -1.3489584e-06, -3.5285944e-07, -9.506044e-05, 6.206637e-05, 8.606192e-06, -1.0958212e-06, -3.5516578e-07, -0.00012474938, 5.6564564e-05, 9.596702e-06, -8.342483e-07, -3.5188424e-07, -0.00015150955, 5.037071e-05, 1.040494e-05, -5.6858164e-07, -3.4325524e-07, -0.00017502453, 4.3604156e-05, 1.1024528e-05, -3.0307976e-07, -3.2959383e-07, -0.00019503887, 3.6389116e-05, 1.1452226e-05, -4.185431e-08, -3.112825e-07, -0.00021135999, 2.8852557e-05, 1.168788e-05, 2.1118834e-07, -2.8876266e-07, -0.00022385905, 2.1122156e-05, 1.1734318e-05, 4.5240088e-07, -2.6252616e-07, -0.00023247086, 1.3324285e-05, 1.1597205e-05, 6.7844275e-07, -2.3310567e-07, -0.0002371926, 5.5821024e-06, 1.1284865e-05, 8.8632163e-07, -2.0106522e-07, -0.00023808192, -1.9862475e-06, 1.080805e-05, 1.0734279e-06, -1.6699035e-07, -0.00023525392, -9.269301e-06, 1.0179707e-05, 1.2375623e-06, -1.3147829e-07, -0.00022887741, -1.6163774e-05, 9.414689e-06, 1.3769558e-06, -9.512833e-08, -0.00021917057, -2.257589e-05, 8.529469e-06, 1.4902831e-06, -5.8532482e-08, -0.00020639582, -2.842251e-05, 7.541826e-06, 1.5766676e-06, -2.226652e-08, -0.0001908543, -3.3632063e-05, 6.4705287e-06, 1.6356801e-06, 1.311837e-08, -0.0001728799, -3.8145266e-05, 5.335007e-06, 1.6673299e-06, 4.7103306e-08, -0.00015283293, -4.191563e-05, 4.155031e-06, 1.6720508e-06, 7.920866e-08, -0.00013109372, -4.4909746e-05, 2.950394e-06, 1.6506789e-06, 1.0900016e-07, -0.00010805603, -4.7107358e-05, 1.7406019e-06, 1.6044269e-06, 1.360941e-07, -8.4120424e-05, -4.8501246e-05, 5.4458303e-07, 1.5348518e-06, 1.6016155e-07, -5.968793e-05, -4.9096885e-05, -6.195867e-07, 1.4438201e-06, 1.8093162e-07, -3.5153746e-05, -4.8911937e-05, -1.734935e-06, 1.3334676e-06, 1.9819372e-07, -1.09013345e-05, -4.797557e-05, -2.7858193e-06, 1.2061573e-06, 2.117987e-07, 1.27031235e-05, -4.6327605e-05, -3.7581237e-06, 1.0644358e-06, 2.2165922e-07, 3.531583e-05, -4.401756e-05, -4.639427e-06, 9.109866e-07, 2.2774888e-07, 5.6619927e-05, -4.1103536e-05, -5.4191373e-06, 7.485846e-07, 2.3010065e-07, 7.632953e-05, -3.7651036e-05, -6.088595e-06, 5.8004986e-07, 2.2880432e-07, 9.419308e-05, -3.37317e-05, -6.6411417e-06, 4.082021e-07, 2.2400322e-07, 0.0001099961, -2.9421984e-05, -7.0721553e-06, 2.3581738e-07, 2.1589014e-07, 0.00012356327, -2.4801822e-05, -7.379054e-06, 6.5586256e-08, 2.0470272e-07, 0.0001347598, -1.9953257e-05, -7.5612647e-06, -9.992489e-08, 1.9071823e-07, 0.00014349222, -1.4959106e-05, -7.6201695e-06, -2.5830948e-07, 1.7424792e-07, 0.00014970833, -9.901651e-06, -7.5590124e-06, -4.0735262e-07, 1.5563107e-07, 0.00015339672, -4.861377e-06, -7.3827896e-06, -5.45059e-07, 1.3522879e-07, 0.00015458548, 8.420873e-08, -7.098112e-06, -6.6967635e-07, 1.1341764e-07, 0.00015334053, 4.861681e-06, -6.7130477e-06, -7.7971447e-07, 9.058333e-08, 0.00014976322, 9.402696e-06, -6.23695e-06, -8.739594e-07, 6.711439e-08, 0.00014398767, 1.364488e-05, -5.680266e-06, -9.514829e-07, 4.339609e-08, 0.00013617745, 1.7532591e-05, -5.05434e-06, -1.0116473e-06, 1.9804533e-08, 0.00012652224, 2.1017559e-05, -4.371206e-06, -1.0541056e-06, -3.2988252e-09, 0.0001152338, 2.4059378e-05, -3.6433796e-06, -1.0787968e-06, -2.5572303e-08, 0.00010254213, 2.662588e-05, -2.8836455e-06, -1.0859374e-06, -4.669862e-08, 8.869116e-05, 2.8693334e-05, -2.1048527e-06, -1.0760084e-06, -6.638898e-08, 7.393456e-05, 3.0246556e-05, -1.3197115e-06, -1.0497396e-06, -8.43866e-08, 5.853149e-05, 3.127883e-05, -5.406018e-07, -1.008089e-06, -1.0046959e-07, 4.274236e-05, 3.1791744e-05, 2.2060745e-07, -9.522209e-07, -1.1445326e-07, 2.6824775e-05, 3.1794883e-05, 9.527252e-07, -8.834806e-07, -1.2619164e-07, 1.1029648e-05, 3.1305397e-05, 1.6453887e-06, -8.0336747e-07, -1.3557855e-07, -4.402484e-06, 3.0347495e-05, 2.2891963e-06, -7.1350655e-07, -1.4254776e-07, -1.9244822e-05, 2.8951832e-05, 2.8758209e-06, -6.156193e-07, -1.4707284e-07, -3.328736e-05, 2.7154802e-05, 3.3981019e-06, -5.114932e-07, -1.4916608e-07, -4.633957e-05, 2.4997797e-05, 3.8501175e-06, -4.0295237e-07, -1.4887705e-07, -5.8232705e-05, 2.2526383e-05, 4.2272345e-06, -2.9182763e-07, -1.4629057e-07, -6.882166e-05, 1.9789464e-05, 4.5261377e-06, -1.7992816e-07, -1.4152423e-07, -7.7986435e-05, 1.6838409e-05, 4.7448334e-06, -6.901412e-08, -1.3472541e-07, -8.563317e-05, 1.3726165e-05, 4.8826405e-06, 3.922905e-08, -1.2606803e-07, -9.169465e-05, 1.0506393e-05, 4.9401533e-06, 1.4321412e-07, -1.15748946e-07, -9.613054e-05, 7.2326084e-06, 4.919189e-06, 2.4147343e-07, -1.0398412e-07, -9.8927005e-05, 3.9573574e-06, 4.8227216e-06, 3.3267753e-07, -9.100465e-08, -0.00010009611, 7.314347e-07, 4.654794e-06, 4.156512e-07, -7.705263e-08, -9.967471e-05, -2.3968441e-06, 4.4204185e-06, 4.8938637e-07, -6.237709e-08, -9.7723074e-05, -5.382307e-06, 4.12547e-06, 5.5305213e-07, -4.722985e-08, -9.432313e-05, -8.18352e-06, 3.7765624e-06, 6.060018e-07, -3.1861553e-08, -8.957648e-05, -1.0763302e-05, 3.3809233e-06, 6.4777635e-07, -1.6517804e-08, -8.360217e-05, -1.3089159e-05, 2.9462597e-06, 6.7810555e-07, -1.4355486e-09, -7.653425e-05, -1.5133629e-05, 2.4806236e-06, 6.969056e-07, 1.316032e-08, -6.851917e-05, -1.6874536e-05, 1.9922754e-06, 7.0427427e-07, 2.7060032e-08, -5.9713133e-05, -1.8295155e-05, 1.489548e-06, 7.00483e-07, 4.0071686e-08, -5.0279305e-05, -1.9384292e-05, 9.807164e-07, 6.859671e-07, 5.2023616e-08, -4.0385075e-05, -2.0136264e-05, 4.738707e-07, 6.6131344e-07, 6.276637e-08, -3.0199322e-05, -2.0550806e-05, -2.320288e-08, 6.2724604e-07, 7.2174274e-08, -1.9889725e-05, -2.063289e-05, -5.031323e-07, 5.8461046e-07, 8.0146584e-08, -9.6202275e-06, -2.039247e-05, -9.5906e-07, 5.343565e-07, 8.66082e-08, 4.5138748e-07, -1.9844165e-05, -1.384732e-06, 4.7751985e-07, 9.1509975e-08, 1.01757305e-05, -1.900687e-05, -1.7745737e-06, 4.1520332e-07, 9.482858e-08, 1.941384e-05, -1.7903314e-05, -2.1237545e-06, 3.4855745e-07, 9.6566005e-08};
endpackage
`endif
