`ifndef COEFFICIENTS_FX_SV_
`define COEFFICIENTS_FX_SV_
package Coefficients_Fx;
	localparam N = 6;
	localparam M = 6;
	localparam COEFF_BIAS = 48;
	localparam logic signed[63:0] Lfr[0:5] = {64'd275737174041358, 64'd275737174041358, 64'd270572062376816, 64'd270572062376816, 64'd267764037443920, 64'd267764037443920};
	localparam logic signed[63:0] Lfi[0:5] = {64'd35027404521307, - 64'd35027404521307, 64'd24610455576128, - 64'd24610455576128, 64'd8786138880886, - 64'd8786138880886};
	localparam logic signed[63:0] Lbr[0:5] = {64'd275737174041358, 64'd275737174041358, 64'd270572062376816, 64'd270572062376816, 64'd267764037443920, 64'd267764037443920};
	localparam logic signed[63:0] Lbi[0:5] = {64'd35027404521307, - 64'd35027404521307, 64'd24610455576128, - 64'd24610455576128, 64'd8786138880886, - 64'd8786138880886};
	localparam logic signed[63:0] Wfr[0:5] = {- 64'd2651298819, - 64'd2651298819, - 64'd1748955530, - 64'd1748955530, - 64'd572084438, - 64'd572084438};
	localparam logic signed[63:0] Wfi[0:5] = {64'd1889252854, - 64'd1889252854, - 64'd672365497, 64'd672365497, - 64'd1400387597, 64'd1400387597};
	localparam logic signed[63:0] Wbr[0:5] = {64'd2651298819, 64'd2651298819, 64'd1748955530, 64'd1748955530, 64'd572084438, 64'd572084438};
	localparam logic signed[63:0] Wbi[0:5] = {- 64'd1889252854, 64'd1889252854, 64'd672365497, - 64'd672365497, 64'd1400387597, - 64'd1400387597};
	localparam logic signed[63:0] Ffr[0:5][0:149] = '{
		'{- 64'd113364990210738416, - 64'd3983886949576016, 64'd5569828753829607, - 64'd257905633687294, - 64'd125531372261044, 64'd19081521365657, - 64'd114421661700765920, - 64'd252787103572623, 64'd5431958010978724, - 64'd364655848560909, - 64'd112480991897162, 64'd20439689021416, - 64'd113632587199134496, 64'd3389547035691944, 64'd5211139927079489, - 64'd462952836698487, - 64'd97966540628453, 64'd21439061241915, - 64'd111056214328367104, 64'd6887404564960130, 64'd4912948569680208, - 64'd551443750702659, - 64'd82255227722555, 64'd22072669137832, - 64'd106777957837526336, 64'd10188757390959440, 64'd4544049735880285, - 64'd628965316574561, - 64'd65626649275951, 64'd22339533300416, - 64'd100908170763820064, 64'd13245995967219460, 64'd4112067807347828, - 64'd694557617108024, - 64'd48368034197952, 64'd22244530428458, - 64'd93579769493015312, 64'd16016576473275068, 64'd3625440673530840, - 64'd747474298852112, - 64'd30769487045376, 64'd21798170151482, - 64'd84945559090488032, 64'd18463571347437996, 64'd3093265326712530, - 64'd787189129275752, - 64'd13119303432000, 64'd21016287831245, - 64'd75175308887683760, 64'd20556116822289656, 64'd2525136816144404, - 64'd813398890629686, 64'd4300569300313, 64'd19919660315895, - 64'd64452631037034520, 64'd22269752907785916, 64'd1930983287264629, - 64'd826022655588578, 64'd21218857579341, 64'd18533552672876, - 64'd52971716570588112, 64'd23586653090378920, 64'd1320899826471287, - 64'd825197546169895, 64'd37379009805054, 64'd16887204824597, - 64'd40933984407312960, 64'd24495742838164032, 64'd704983783260547, - 64'd811271130823059, 64'd52542909780549, 64'd15013267744604, - 64'd28544698759471100, 64'd24992707792833616, 64'd93174151604766, - 64'd784790664188415, 64'd66494204647644, 64'd12947199433882, - 64'd16009609512006336, 64'd25079894261453868, - 64'd504902536308573, - 64'd746489419146093, 64'd79041203994704, 64'd10726631282315, - 64'd3531668426439428, 64'd24766106268687644, - 64'd1080077515416534, - 64'd697270400804040, 64'd90019314700874, 64'd8390715627535, 64'd8692128499272152, 64'd24066304968969788, - 64'd1623774200497883, - 64'd638187766502393, 64'd99292984344543, 64'd5979465353495, 64'd20473725441161716, 64'd23001217626535588, - 64'd2128129839791589, - 64'd570426304329795, 64'd106757134494146, 64'd3533096228055, 64'd31636774781455288, 64'd21596864629957068, - 64'd2586102792344198, - 64'd495279344753834, 64'd112338073775578, 64'd1091382369241, 64'd42019150127781576, 64'd19884014100661044, - 64'd2991564080733010, - 64'd414125495567832, 64'd115993889134106, - 64'd1306965237301, 64'd51475170700469208, 64'd17897574568536412, - 64'd3339372154386992, - 64'd328404599363619, 64'd117714322045471, - 64'd3624887860422, 64'd59877508894710776, 64'd15675936912113984, - 64'd3625430092182028, - 64'd239593315175250, 64'd117520144452945, - 64'd5827527222024, 64'd67118758563459712, 64'd13260277289108012, - 64'd3846724771409130, - 64'd149180721926746, 64'd115462056794691, - 64'd7882725072588, 64'd73112647520344288, 64'd10693833111819658, - 64'd4001347828734964, - 64'd58644331081793, 64'd111619137529093, - 64'd9761467408887, 64'd77794883829637216, 64'd8021164250755380, - 64'd4088498532644028, 64'd30573120247393, 64'd106096879966224, - 64'd11438267646808, 64'd81123631533078432, 64'd5287411581728942, - 64'd4108468971513664, 64'd117085746117695, 64'd99024857885551, - 64'd12891484174376},
		'{- 64'd113364990210668768, - 64'd3983886949580926, 64'd5569828753831866, - 64'd257905633687862, - 64'd125531372260965, 64'd19081521365658, - 64'd114421661700723616, - 64'd252787103575427, 64'd5431958010980114, - 64'd364655848561268, - 64'd112480991897113, 64'd20439689021417, - 64'd113632587199119552, 64'd3389547035691238, 64'd5211139927080010, - 64'd462952836698636, - 64'd97966540628433, 64'd21439061241916, - 64'd111056214328379040, 64'd6887404564961484, 64'd4912948569679872, - 64'd551443750702600, - 64'd82255227722564, 64'd22072669137833, - 64'd106777957837564336, 64'd10188757390962776, 64'd4544049735879120, - 64'd628965316574301, - 64'd65626649275989, 64'd22339533300417, - 64'd100908170763882864, 64'd13245995967224680, 64'd4112067807345872, - 64'd694557617107572, - 64'd48368034198017, 64'd22244530428459, - 64'd93579769493101280, 64'd16016576473282042, 64'd3625440673528145, - 64'd747474298851480, - 64'd30769487045467, 64'd21798170151483, - 64'd84945559090595232, 64'd18463571347446564, 64'd3093265326709158, - 64'd787189129274954, - 64'd13119303432114, 64'd21016287831246, - 64'd75175308887809968, 64'd20556116822299648, 64'd2525136816140422, - 64'd813398890628739, 64'd4300569300178, 64'd19919660315896, - 64'd64452631037177248, 64'd22269752907797136, 64'd1930983287260118, - 64'd826022655587501, 64'd21218857579189, 64'd18533552672878, - 64'd52971716570744688, 64'd23586653090391160, 64'd1320899826466332, - 64'd825197546168708, 64'd37379009804886, 64'd16887204824598, - 64'd40933984407480536, 64'd24495742838177072, 64'd704983783255237, - 64'd811271130821784, 64'd52542909780369, 64'd15013267744605, - 64'd28544698759646752, 64'd24992707792847228, 64'd93174151599195, - 64'd784790664187074, 64'd66494204647454, 64'd12947199433883, - 64'd16009609512187064, 64'd25079894261467816, - 64'd504902536314311, - 64'd746489419144709, 64'd79041203994508, 64'd10726631282316, - 64'd3531668426622232, 64'd24766106268701704, - 64'd1080077515422342, - 64'd697270400802637, 64'd90019314700676, 64'd8390715627536, 64'd8692128499090228, 64'd24066304968983732, - 64'd1623774200503669, - 64'd638187766500992, 64'd99292984344346, 64'd5979465353495, 64'd20473725440983556, 64'd23001217626549200, - 64'd2128129839797260, - 64'd570426304328420, 64'd106757134493953, 64'd3533096228056, 64'd31636774781283612, 64'd21596864629970132, - 64'd2586102792349668, - 64'd495279344752505, 64'd112338073775392, 64'd1091382369241, 64'd42019150127618968, 64'd19884014100673372, - 64'd2991564080738195, - 64'd414125495566571, 64'd115993889133928, - 64'd1306965237301, 64'd51475170700318016, 64'd17897574568547828, - 64'd3339372154391818, - 64'd328404599362442, 64'd117714322045306, - 64'd3624887860422, 64'd59877508894573136, 64'd15675936912124328, - 64'd3625430092186428, - 64'd239593315174175, 64'd117520144452794, - 64'd5827527222024, 64'd67118758563337464, 64'd13260277289117144, - 64'd3846724771413042, - 64'd149180721925787, 64'd115462056794557, - 64'd7882725072588, 64'd73112647520238992, 64'd10693833111827464, - 64'd4001347828738340, - 64'd58644331080962, 64'd111619137528977, - 64'd9761467408887, 64'd77794883829550112, 64'd8021164250761770, - 64'd4088498532646828, 64'd30573120248085, 64'd106096879966127, - 64'd11438267646808, 64'd81123631533010496, 64'd5287411581733847, - 64'd4108468971515856, 64'd117085746118241, 64'd99024857885475, - 64'd12891484174376},
		'{- 64'd261185979523892064, - 64'd22456890558529396, 64'd8607393505184881, - 64'd1769784954461006, 64'd241447559502841, 64'd1933593015434, - 64'd270800817222180096, - 64'd16047694531985916, 64'd7900070649760353, - 64'd1716378903106676, 64'd254857519535561, - 64'd3773288418972, - 64'd277282227462791680, - 64'd9929647949627100, 64'd7168828679240094, - 64'd1650925382366498, 64'd265020553967774, - 64'd9055741381813, - 64'd280785027968515808, - 64'd4138808128063452, 64'd6421989129967633, - 64'd1574846110810426, 64'd272065566502174, - 64'd13894456389570, - 64'd281480698205836832, 64'd1294223557194100, 64'd5667447612258315, - 64'd1489562841760350, 64'd276141168090658, - 64'd18275501295111, - 64'd279554672781074240, 64'd6344208747836490, 64'd4912630705697034, - 64'd1396484358864565, 64'd277412971381418, - 64'd22190081292982, - 64'd275203692143743456, 64'd10991136482630424, 64'd4164460088880028, - 64'd1296994478805553, 64'd276060914540424, - 64'd25634268340864, - 64'd268633230909669152, 64'd15220049038531744, 64'd3429323737345382, - 64'd1192441102045094, 64'd272276636914191, - 64'd28608704561309, - 64'd260055022018696416, 64'd19020833458887984, 64'd2713053970157080, - 64'd1084126340131656, 64'd266260926991562, - 64'd31118284113950, - 64'd249684692820901536, 64'd22387983019644088, 64'd2020912077975607, - 64'd973297736300737, 64'd258221261063288, - 64'd33171817918496, - 64'd237739527061999296, 64'd25320332868942032, 64'd1357579223514040, - 64'd861140584957512, 64'd248369448891663, - 64'd34781685466361, - 64'd224436364632737920, 64'd27820774022308884, 64'd727153269036316, - 64'd748771345199828, 64'd236919400609314, - 64'd35963477787308, - 64'd209989648876552352, 64'd29895949807821008, 64'd133151154946584, - 64'd637232133865376, 64'd224085026986094, - 64'd36735635440535, - 64'd194609629231121920, 64'd31555938736379624, - 64'd421483571559838, - 64'd527486274706295, 64'd210078283153949, - 64'd37119085180767, - 64'd178500725027667200, 64'd32813927624776528, - 64'd934368498510874, - 64'd420414872234720, 64'd195107363878338, - 64'd37136878712585, - 64'd161860054400109248, 64'd33685878626842608, - 64'd1403665797068552, - 64'd316814371561296, 64'd179375056526202, - 64'd36813836693955, - 64'd144876130476242112, 64'd34190193633935372, - 64'd1828061820100178, - 64'd217395059174395, 64'd163077256018137, - 64'd36176200885914, - 64'd127727725344849952, 64'd34347379293590144, - 64'd2206743300987920, - 64'd122780454080956, 64'd146401644278134, - 64'd35251297072942, - 64'd110582900724628400, 64'd34179715667531056, - 64'd2539370602628581, - 64'd33507534043250, 64'd129526535018160, - 64'd34067211100752, - 64'd93598202809657440, 64'd33710931310532892, - 64'd2826048462808806, 64'd49972262215125, 64'd112619883125651, - 64'd32652480097898, - 64'd76918017437303328, 64'd32965887302861392, - 64'd3067294674551256, 64'd127291319017218, 64'd95838456466683, - 64'd31035800667583, - 64'd60674080521596304, 64'd31970272514089748, - 64'd3264007128945235, 64'd198163478416821, 64'd79327166581764, - 64'd29245755558798, - 64'd44985137620731944, 64'd30750312117747640, - 64'd3417429633740691, 64'd262381091554607, 64'd63218553538739, - 64'd27310560053785, - 64'd29956745562421616, 64'd29332491117099896, - 64'd3529116903943056, 64'd319811553507675, 64'd47632419121166, - 64'd25257829044054, - 64'd15681208235173768, 64'd27743294384802212, - 64'd3600899101145688, 64'd370393388611762, 64'd32675601571658, - 64'd23114365511491},
		'{- 64'd261185979523428576, - 64'd22456890558562344, 64'd8607393505199444, - 64'd1769784954464604, 64'd241447559503349, 64'd1933593015434, - 64'd270800817221775808, - 64'd16047694532014440, 64'd7900070649773052, - 64'd1716378903109822, 64'd254857519536005, - 64'd3773288418972, - 64'd277282227462446208, - 64'd9929647949651234, 64'd7168828679250940, - 64'd1650925382369192, 64'd265020553968155, - 64'd9055741381813, - 64'd280785027968228288, - 64'd4138808128083280, 64'd6421989129976653, - 64'd1574846110812677, 64'd272065566502491, - 64'd13894456389570, - 64'd281480698205605952, 64'd1294223557178464, 64'd5667447612265551, - 64'd1489562841762165, 64'd276141168090914, - 64'd18275501295111, - 64'd279554672780898240, 64'd6344208747824902, 64'd4912630705702542, - 64'd1396484358865959, 64'd277412971381615, - 64'd22190081292981, - 64'd275203692143620224, 64'd10991136482622716, 64'd4164460088883876, - 64'd1296994478806542, 64'd276060914540563, - 64'd25634268340863, - 64'd268633230909596192, 64'd15220049038527722, 64'd3429323737347648, - 64'd1192441102045696, 64'd272276636914275, - 64'd28608704561307, - 64'd260055022018670912, 64'd19020833458887424, 64'd2713053970157851, - 64'd1084126340131892, 64'd266260926991594, - 64'd31118284113949, - 64'd249684692820920544, 64'd22387983019646772, 64'd2020912077974979, - 64'd973297736300630, 64'd258221261063272, - 64'd33171817918495, - 64'd237739527062059552, 64'd25320332868947704, 64'd1357579223512113, - 64'd861140584957086, 64'd248369448891602, - 64'd34781685466359, - 64'd224436364632836096, 64'd27820774022317292, 64'd727153269033198, - 64'd748771345199110, 64'd236919400609212, - 64'd35963477787306, - 64'd209989648876684928, 64'd29895949807831892, 64'd133151154942383, - 64'd637232133864391, 64'd224085026985954, - 64'd36735635440533, - 64'd194609629231285376, 64'd31555938736392708, - 64'd421483571565008, - 64'd527486274705071, 64'd210078283153775, - 64'd37119085180765, - 64'd178500725027857888, 64'd32813927624791544, - 64'd934368498516900, - 64'd420414872233284, 64'd195107363878135, - 64'd37136878712583, - 64'd161860054400323584, 64'd33685878626859292, - 64'd1403665797075320, - 64'd316814371559676, 64'd179375056525972, - 64'd36813836693953, - 64'd144876130476476512, 64'd34190193633953452, - 64'd1828061820107576, - 64'd217395059172618, 64'd163077256017885, - 64'd36176200885912, - 64'd127727725345100896, 64'd34347379293609364, - 64'd2206743300995836, - 64'd122780454079049, 64'd146401644277863, - 64'd35251297072941, - 64'd110582900724892480, 64'd34179715667551152, - 64'd2539370602636909, - 64'd33507534041241, 64'd129526535017876, - 64'd34067211100751, - 64'd93598202809931344, 64'd33710931310553636, - 64'd2826048462817442, 64'd49972262217212, 64'd112619883125355, - 64'd32652480097896, - 64'd76918017437583840, 64'd32965887302882540, - 64'd3067294674560098, 64'd127291319019360, 64'd95838456466380, - 64'd31035800667582, - 64'd60674080521880440, 64'd31970272514111080, - 64'd3264007128954190, 64'd198163478418993, 64'd79327166581456, - 64'd29245755558796, - 64'd44985137621016856, 64'd30750312117768944, - 64'd3417429633749668, 64'd262381091556787, 64'd63218553538431, - 64'd27310560053784, - 64'd29956745562704656, 64'd29332491117120984, - 64'd3529116903951972, 64'd319811553509842, 64'd47632419120859, - 64'd25257829044053, - 64'd15681208235452464, 64'd27743294384822912, - 64'd3600899101154465, 64'd370393388613898, 64'd32675601571355, - 64'd23114365511490},
		'{- 64'd147927123522367456, - 64'd18177492446279264, 64'd3137698184896970, - 64'd1488192028122724, 64'd338884941609365, - 64'd83132750190217, - 64'd156324607661916704, - 64'd15447556199019812, 64'd2572490864587542, - 64'd1349781309511470, 64'd311842990457516, - 64'd77626660430557, - 64'd163408861711848480, - 64'd12922733796088518, 64'd2051844969362986, - 64'd1219873695525226, 64'd286301234270640, - 64'd72378730192471, - 64'd169279715903773056, - 64'd10592180041143310, 64'd1573311048560416, - 64'd1098104073152683, 64'd262204033560234, - 64'd67382238575553, - 64'd174031670337643904, - 64'd8445419759004248, 64'd1134529129707866, - 64'd984114438549139, 64'd239496148021515, - 64'd62630255352860, - 64'd177754080110616032, - 64'd6472348047584440, 64'd733228199975529, - 64'd877554426523398, 64'd218122883876100, - 64'd58115683859598, - 64'd180531340250850880, - 64'd4663229266772438, 64'd367225438650931, - 64'd778081764645723, 64'd198030225524146, - 64'd53831300404132, - 64'd182443069855621344, - 64'd3008694886471708, 64'd34425226629464, - 64'd685362657548161, 64'd179164952541371, - 64'd49769790396593, - 64'd183564294892240736, - 64'd1499740308324762, - 64'd267182042787098, - 64'd599072106698097, 64'd161474743008033, - 64'd45923781382925, - 64'd183965629175753376, - 64'd127720768310654, - 64'd539521329111766, - 64'd518894170645069, 64'd144908264109849, - 64'd42285873164940, - 64'd183713453089154848, 64'd1115653579602926, - 64'd784434464784578, - 64'd444522170469735, 64'd129415250904971, - 64'd38848665179692, - 64'd182870089660314496, 64'd2238323305255050, - 64'd1003681810516536, - 64'd375658844902448, 64'd114946574106669, - 64'd35604781304352, - 64'd181493977654918944, 64'd3247885982404254, - 64'd1198944027602716, - 64'd312016459327057, 64'd101454297688191, - 64'd32546892245770, - 64'd179639841386790816, 64'd4151603026088577, - 64'd1371823950268495, - 64'd253316872643342, 64'd88891727074462, - 64'd29667735666990, - 64'd177358856986020544, 64'd4956407011924468, - 64'd1523848542371368, - 64'd199291565728716, 64'd77213448644859, - 64'd26960134196258, - 64'd174698814901622912, 64'd5668909407507587, - 64'd1656470923973247, - 64'd149681635016508, 64'd66375361232269, - 64'd24417011457433, - 64'd171704278449040032, 64'd6295408651269154, - 64'd1771072454427026, - 64'd104237754493935, 64'd56334700265924, - 64'd22031406254313, - 64'd168416738243893632, 64'd6841898519060024, - 64'd1868964859688488, - 64'd62720109217924, 64'd47050055169258, - 64'd19796485035030, - 64'd164874762392079616, 64'd7314076723390628, - 64'd1951392392572694, - 64'd24898303250727, 64'd38481380589084, - 64'd17705552756628, - 64'd161114142332723552, 64'd7717353694656953, - 64'd2019534015624960, 64'd9448755270026, 64'd30590001998816, - 64'd15752062263952, - 64'd157168034254798720, 64'd8056861497840441, - 64'd2074505597172628, 64'd40532989391103, 64'd23338616186249, - 64'd13929622291208, - 64'd153067096030477760, 64'd8337462842091858, - 64'd2117362111967220, 64'd68557306567997, 64'd16691287105506, - 64'd12232004189014, - 64'd148839619628647360, 64'd8563760144304924, - 64'd2149099838619291, 64'd93715767650942, 64'd10613437543130, - 64'd10653147474290, - 64'd144511658990586496, 64'd8740104611263724, - 64'd2170658546772659, 64'd116193769584212, 64'd5071837020033, - 64'd9187164295181, - 64'd140107153366689824, 64'd8870605308217606, - 64'd2182923667662533, 64'd136168239917123, 64'd34586323870, - 64'd7828342898123},
		'{- 64'd147927123521392000, - 64'd18177492446348480, 64'd3137698184927293, - 64'd1488192028130171, 64'd338884941610422, - 64'd83132750190221, - 64'd156324607660996992, - 64'd15447556199085032, 64'd2572490864616129, - 64'd1349781309518492, 64'd311842990458513, - 64'd77626660430561, - 64'd163408861710982336, - 64'd12922733796149900, 64'd2051844969389905, - 64'd1219873695531840, 64'd286301234271579, - 64'd72378730192475, - 64'd169279715902958368, - 64'd10592180041201008, 64'd1573311048585734, - 64'd1098104073158904, 64'd262204033561118, - 64'd67382238575556, - 64'd174031670336878528, - 64'd8445419759058417, 64'd1134529129731650, - 64'd984114438554984, 64'd239496148022345, - 64'd62630255352863, - 64'd177754080109897920, - 64'd6472348047635232, 64'd733228199997842, - 64'd877554426528883, 64'd218122883876879, - 64'd58115683859601, - 64'd180531340250177952, - 64'd4663229266820000, 64'd367225438671837, - 64'd778081764650863, 64'd198030225524876, - 64'd53831300404135, - 64'd182443069854991616, - 64'd3008694886516184, 64'd34425226649026, - 64'd685362657552972, 64'd179164952542054, - 64'd49769790396595, - 64'd183564294891652288, - 64'd1499740308366294, - 64'd267182042768819, - 64'd599072106702593, 64'd161474743008671, - 64'd45923781382927, - 64'd183965629175204256, - 64'd127720768349380, - 64'd539521329094712, - 64'd518894170649265, 64'd144908264110445, - 64'd42285873164942, - 64'd183713453088643200, 64'd1115653579566872, - 64'd784434464768689, - 64'd444522170473645, 64'd129415250905526, - 64'd38848665179694, - 64'd182870089659838528, 64'd2238323305221536, - 64'd1003681810501757, - 64'd375658844906086, 64'd114946574107185, - 64'd35604781304353, - 64'd181493977654476864, 64'd3247885982373158, - 64'd1198944027588991, - 64'd312016459330436, 64'd101454297688671, - 64'd32546892245771, - 64'd179639841386380928, 64'd4151603026059772, - 64'd1371823950255771, - 64'd253316872646475, 64'd88891727074907, - 64'd29667735666992, - 64'd177358856985641184, 64'd4956407011897833, - 64'd1523848542359593, - 64'd199291565731617, 64'd77213448645271, - 64'd26960134196259, - 64'd174698814901272480, 64'd5668909407483011, - 64'd1656470923962372, - 64'd149681635019187, 64'd66375361232649, - 64'd24417011457435, - 64'd171704278448716992, 64'd6295408651246523, - 64'd1771072454417002, - 64'd104237754496406, 64'd56334700266274, - 64'd22031406254314, - 64'd168416738243596480, 64'd6841898519039232, - 64'd1868964859679269, - 64'd62720109220197, 64'd47050055169581, - 64'd19796485035031, - 64'd164874762391806912, 64'd7314076723371573, - 64'd1951392392564236, - 64'd24898303252813, 64'd38481380589380, - 64'd17705552756629, - 64'd161114142332473920, 64'd7717353694639534, - 64'd2019534015617218, 64'd9448755268116, 64'd30590001999087, - 64'd15752062263952, - 64'd157168034254570816, 64'd8056861497824561, - 64'd2074505597165561, 64'd40532989389359, 64'd23338616186497, - 64'd13929622291209, - 64'd153067096030270272, 64'd8337462842077426, - 64'd2117362111960788, 64'd68557306566409, 64'd16691287105731, - 64'd12232004189015, - 64'd148839619628459104, 64'd8563760144291853, - 64'd2149099838613457, 64'd93715767649500, 64'd10613437543335, - 64'd10653147474290, - 64'd144511658990416288, 64'd8740104611251929, - 64'd2170658546767385, 64'd116193769582909, 64'd5071837020218, - 64'd9187164295182, - 64'd140107153366536528, 64'd8870605308207004, - 64'd2182923667657784, 64'd136168239915949, 64'd34586324037, - 64'd7828342898124}};
	localparam logic signed[63:0] Ffi[0:5][0:149] = '{
		'{64'd27061454864742516, - 64'd29329963185269764, 64'd195520791088329, 64'd900075992202870, - 64'd84307738655099, - 64'd14039756020202, 64'd12402408768204324, - 64'd29227842841782012, 64'd884657663660782, 64'd849633769750120, - 64'd98210562395013, - 64'd11379009668686, - 64'd2089310716763816, - 64'd28663497405476736, 64'd1542589681822757, 64'd786935553955462, - 64'd110205960410614, - 64'd8603488459578, - 64'd16187425555932316, - 64'd27657395440758048, 64'd2159630788206751, 64'd713283119733266, - 64'd120150622728524, - 64'd5760181395202, - 64'd29677543699628088, - 64'd26236521060170792, 64'd2726986023501624, 64'd630120057110324, - 64'd127937412862532, - 64'd2895986842769, - 64'd42360272641980240, - 64'd24433782808960836, 64'd3236869219002734, 64'd539005289400233, - 64'd133496171871328, - 64'd56969036973, - 64'd54054017037580968, - 64'd22287343042577064, 64'd3682601721153442, 64'd441585415965900, - 64'd136793914424840, 64'd2712353664127, - 64'd64597423746336640, - 64'd19839880438164920, 64'd4058691049914580, 64'd339566348590174, - 64'd137834428881022, 64'd5369678241846, - 64'd73851444194581232, - 64'd17137799030007612, 64'd4360888739188662, 64'd234684710043639, - 64'd136657302553573, 64'd7875534604264, - 64'd81700990774571280, - 64'd14230397676234388, 64'd4586226957255934, 64'd128679455567068, - 64'd133336401964652, 64'd10193842767793, - 64'd88056171038730048, - 64'd11169014147466116, 64'd4733033852605743, 64'd23264162984228, - 64'd127977845802236, 64'd12292402275104, - 64'd92853090562627088, - 64'd8006158078720994, 64'd4800927910201560, - 64'd79899584555584, - 64'd120717515430476, 64'd14143307752129, - 64'd96054222436410784, - 64'd4794646848838514, 64'd4790791929893918, - 64'd179227327124325, - 64'd111718154039706, 64'd15723285832956, - 64'd97648348286379680, - 64'd1586758055376818, 64'd4704727547520385, - 64'd273235005292775, - 64'd101166110793507, 64'd17013950050470, - 64'd97650082419767936, 64'd1566588350849615, 64'd4545991505738860, - 64'd360560062034348, - 64'd89267790573839, 64'd18001971679645, - 64'd96098997026461056, 64'd4616606003936770, 64'd4318915141828897, - 64'd439980087802016, - 64'd76245873099580, 64'd18679165906927, - 64'd93058372269148240, 64'd7517364837884810, 64'd4028808790082756, - 64'd510428773391513, - 64'd62335367275175, 64'd19042494061181, - 64'd88613600465584832, 64'd10226450409772886, 64'd3681852994070874, - 64'd571008983867665, - 64'd47779567608419, 64'd19093983958108, - 64'd82870278340830400, 64'd12705550923365190, 64'd3284978586676226, - 64'd621002817253347, - 64'd32825979431485, 64'd18840571661139, - 64'd75952025442497056, 64'd14920964416583992, 64'd2845737821634594, - 64'd659878563016750, - 64'd17722278495844, 64'd18293869129252, - 64'd67998070219142936, 64'd16844020033214614, 64'd2372168828306202, - 64'd687294526803150, - 64'd2712368334485, 64'd17469863289503, - 64'd59160647924404656, 64'd18451408816580252, 64'd1872655711080900, - 64'd703099738523027, 64'd11967404346242, 64'd16388553024781, - 64'd49602256403463392, 64'd19725421015109816, 64'd1355786626346778, - 64'd707331610041940, 64'd26091819994366, 64'd15073531393143, - 64'd39492816932973920, 64'd20654088451171928, 64'd830212144096177, - 64'd700210655575872, 64'd39450090815028, 64'd13551521084012, - 64'd29006787622315340, 64'd21231232050203092, 64'd304506139344359, - 64'd682132431790285, 64'd51848853708365, 64'd11851871661078},
		'{- 64'd27061454864950924, 64'd29329963185285884, - 64'd195520791094942, - 64'd900075992201277, 64'd84307738654874, 64'd14039756020203, - 64'd12402408768417152, 64'd29227842841798412, - 64'd884657663667541, - 64'd849633769748489, 64'd98210562394782, 64'd11379009668687, 64'd2089310716550064, 64'd28663497405493156, - 64'd1542589681829552, - 64'd786935553953819, 64'd110205960410382, 64'd8603488459578, 64'd16187425555721056, 64'd27657395440774216, - 64'd2159630788213471, - 64'd713283119731638, 64'd120150622728295, 64'd5760181395203, 64'd29677543699422628, 64'd26236521060186464, - 64'd2726986023508166, - 64'd630120057108737, 64'd127937412862309, 64'd2895986842770, 64'd42360272641783696, 64'd24433782808975776, - 64'd3236869219008998, - 64'd539005289398711, 64'd133496171871114, 64'd56969036974, 64'd54054017037396248, 64'd22287343042591052, - 64'd3682601721159334, - 64'd441585415964465, 64'd136793914424639, - 64'd2712353664127, 64'd64597423746166368, 64'd19839880438177752, - 64'd4058691049920017, - 64'd339566348588847, 64'd137834428880836, - 64'd5369678241846, 64'd73851444194427808, 64'd17137799030019116, - 64'd4360888739193568, - 64'd234684710042438, 64'd136657302553405, - 64'd7875534604264, 64'd81700990774436672, 64'd14230397676244412, - 64'd4586226957260245, - 64'd128679455566009, 64'd133336401964504, - 64'd10193842767793, 64'd88056171038615952, 64'd11169014147474542, - 64'd4733033852609405, - 64'd23264162983325, 64'd127977845802110, - 64'd12292402275104, 64'd92853090562534800, 64'd8006158078727724, - 64'd4800927910204531, 64'd79899584556320, 64'd120717515430374, - 64'd14143307752129, 64'd96054222436341232, 64'd4794646848843485, - 64'd4790791929896167, 64'd179227327124888, 64'd111718154039628, - 64'd15723285832956, 64'd97648348286333408, 64'd1586758055379994, - 64'd4704727547521895, 64'd273235005293160, 64'd101166110793454, - 64'd17013950050471, 64'd97650082419745088, - 64'd1566588350848240, - 64'd4545991505739625, 64'd360560062034553, 64'd89267790573811, - 64'd18001971679646, 64'd96098997026461440, - 64'd4616606003937172, - 64'd4318915141828924, 64'd439980087802041, 64'd76245873099577, - 64'd18679165906928, 64'd93058372269171232, - 64'd7517364837886940, - 64'd4028808790082064, 64'd510428773391364, 64'd62335367275197, - 64'd19042494061182, 64'd88613600465629536, - 64'd10226450409776666, - 64'd3681852994069489, 64'd571008983867348, 64'd47779567608464, - 64'd19093983958110, 64'd82870278340895552, - 64'd12705550923370520, - 64'd3284978586674188, 64'd621002817252871, 64'd32825979431553, - 64'd18840571661141, 64'd75952025442581120, - 64'd14920964416590748, - 64'd2845737821631954, 64'd659878563016127, 64'd17722278495933, - 64'd18293869129253, 64'd67998070219244096, - 64'd16844020033222652, - 64'd2372168828303015, 64'd687294526802393, 64'd2712368334593, - 64'd17469863289504, 64'd59160647924520880, - 64'd18451408816589412, - 64'd1872655711077230, 64'd703099738522152, - 64'd11967404346118, - 64'd16388553024782, 64'd49602256403592464, - 64'd19725421015119928, - 64'd1355786626342696, 64'd707331610040964, - 64'd26091819994228, - 64'd15073531393144, 64'd39492816933113472, - 64'd20654088451182804, - 64'd830212144091758, 64'd700210655574812, - 64'd39450090814878, - 64'd13551521084013, 64'd29006787622462876, - 64'd21231232050214544, - 64'd304506139339682, 64'd682132431789160, - 64'd51848853708206, - 64'd11851871661079},
		'{64'd225677438598042560, - 64'd63354485394154200, 64'd4276556762928860, 64'd173233147734769, - 64'd260338546982839, 64'd64414188308395, 64'd194099328777530528, - 64'd62863947226030400, 64'd4863482625348990, 64'd11783768817828, - 64'd229143648540106, 64'd62088170629478, 64'd162903732143129920, - 64'd61832029002577360, 64'd5365829956533783, - 64'd138742379771980, - 64'd197984597261583, 64'd59353276176248, 64'd132349799862027520, - 64'd60305157375926432, 64'd5784783558645604, - 64'd277715051368705, - 64'd167143895985067, 64'd56262452200578, 64'd102673108580712048, - 64'd58331113296847152, 64'd6122209925009098, - 64'd404652718271066, - 64'd136881834266162, 64'd52868283349588, 64'd74085116781183136, - 64'd55958502521860016, 64'd6380593594475096, - 64'd519216814161826, - 64'd107435625726572, 64'd49222535549607, 64'd46772878844103376, - 64'd53236254754919808, 64'd6562972202281639, - 64'd621205062519008, - 64'd79018815374206, 64'd45375738541443, 64'd20899001826037872, - 64'd50213154047608856, 64'd6672870910438875, - 64'd710544014480569, - 64'd51820943869420, 64'd41376808243854, - 64'd3398171237329920, - 64'd46937402616638520, 64'd6714236859671300, - 64'd787280918418317, - 64'd26007454251939, 64'd37272709677485, - 64'd26004168655667776, - 64'd43456219784353120, 64'd6691374240886772, - 64'd851575041235286, - 64'd1719825415355, 64'd33108160760582, - 64'd46827805932517792, - 64'd39815477310187040, 64'd6608880537620060, - 64'd903688558214912, 64'd20924084383897, 64'd28925376892742, - 64'd65800428562538304, - 64'd36059371961594712, 64'd6471584442512415, - 64'd943977124213681, 64'd41829501475068, 64'd24763855875645, - 64'd82875000525838496, - 64'd32230135774440352, 64'd6284485901207953, - 64'd972880234196613, 64'd60924026236796, 64'd20660202381705, - 64'd98025057357911808, - 64'd28367784077415996, 64'd6052698686615020, - 64'd990911475662388, 64'd78156766495518, 64'd16647990873758, - 64'd111243542622272928, - 64'd24509901004605992, 64'd5781395855809029, - 64'd998648769487086, 64'd93497333446865, 64'd12757665602248, - 64'd122541546392837312, - 64'd20691461896333824, 64'd5475758391422012, - 64'd996724689226150, 64'd106934718675527, 64'd9016476061142, - 64'd131946963977888080, - 64'd16944691692066244, 64'd5140927279618252, - 64'd985816942044687, 64'd118476070667219, 64'd5448446070101, - 64'd139503092601186624, - 64'd13298958151233642, 64'd4781959228102836, - 64'd966639087285579, 64'd128145388868866, 64'd2074374468180, - 64'd145267183112758496, - 64'd9780698498861298, 64'd4403786180421141, - 64'd939931561318297, 64'd135982152873408, - 64'd1088134747168, - 64'd149308963046665856, - 64'd6413377883100207, 64'd4011178737413532, - 64'd906453069820362, 64'd142039903698047, - 64'd4024615123238, - 64'd151709146490235968, - 64'd3217477851025686, 64'd3608713553383575, - 64'd866972401104986, 64'd146384793403475, - 64'd6723655676905, - 64'd152557945293218496, - 64'd210512897101834, 64'd3200744733573030, - 64'd822260706594790, 64'd149094118481018, - 64'd9176796484705, - 64'd151953595140436224, 64'd2592926985084004, 64'd2791379221127652, - 64'd773084287119666, 64'd150254851529052, - 64'd11378404419024, - 64'd150000908951570592, 64'd5181109913623697, 64'd2384456126060925, - 64'd720197916448334, 64'd149962184763518, - 64'd13325531523291, - 64'd146809868970240064, 64'd7545074127451866, 64'd1983529915917913, - 64'd664338726404090, 64'd148318097873680, - 64'd15017758507562},
		'{- 64'd225677438598514048, 64'd63354485394190232, - 64'd4276556762943734, - 64'd173233147731185, 64'd260338546982331, - 64'd64414188308392, - 64'd194099328778024256, 64'd62863947226067920, - 64'd4863482625364560, - 64'd11783768814068, 64'd229143648539574, - 64'd62088170629475, - 64'd162903732143639872, 64'd61832029002615920, - 64'd5365829956549861, 64'd138742379775869, 64'd197984597261032, - 64'd59353276176245, - 64'd132349799862547968, 64'd60305157375965608, - 64'd5784783558662007, 64'd277715051372679, 64'd167143895984504, - 64'd56262452200575, - 64'd102673108581237456, 64'd58331113296886536, - 64'd6122209925025654, 64'd404652718275083, 64'd136881834265593, - 64'd52868283349585, - 64'd74085116781708352, 64'd55958502521899248, - 64'd6380593594491644, 64'd519216814165847, 64'd107435625726003, - 64'd49222535549604, - 64'd46772878844623648, 64'd53236254754958536, - 64'd6562972202298028, 64'd621205062522994, 64'd79018815373642, - 64'd45375738541441, - 64'd20899001826548768, 64'd50213154047646760, - 64'd6672870910454965, 64'd710544014484487, 64'd51820943868866, - 64'd41376808243852, 64'd3398171236832432, 64'd46937402616675296, - 64'd6714236859686965, 64'd787280918422136, 64'd26007454251399, - 64'd37272709677482, 64'd26004168655187328, 64'd43456219784388528, - 64'd6691374240901898, 64'd851575041238978, 64'd1719825414833, - 64'd33108160760581, 64'd46827805932057600, 64'd39815477310220848, - 64'd6608880537634544, 64'd903688558218452, - 64'd20924084384398, - 64'd28925376892740, 64'd65800428562101232, 64'd36059371961626704, - 64'd6471584442526171, 64'd943977124217046, - 64'd41829501475544, - 64'd24763855875643, 64'd82875000525426944, 64'd32230135774470372, - 64'd6284485901220903, 64'd972880234199785, - 64'd60924026237245, - 64'd20660202381703, 64'd98025057357527776, 64'd28367784077443900, - 64'd6052698686627101, 64'd990911475665351, - 64'd78156766495936, - 64'd16647990873756, 64'd111243542621918048, 64'd24509901004631672, - 64'd5781395855820190, 64'd998648769489827, - 64'd93497333447253, - 64'd12757665602247, 64'd122541546392512864, 64'd20691461896357200, - 64'd5475758391432213, 64'd996724689228659, - 64'd106934718675882, - 64'd9016476061141, 64'd131946963977594928, 64'd16944691692087254, - 64'd5140927279627466, 64'd985816942046958, - 64'd118476070667540, - 64'd5448446070100, 64'd139503092600925328, 64'd13298958151252256, - 64'd4781959228111047, 64'd966639087287606, - 64'd128145388869152, - 64'd2074374468179, 64'd145267183112529280, 64'd9780698498877512, - 64'd4403786180428342, 64'd939931561320079, - 64'd135982152873659, 64'd1088134747169, 64'd149308963046468608, 64'd6413377883114036, - 64'd4011178737419725, 64'd906453069821900, - 64'd142039903698264, 64'd4024615123238, 64'd151709146490070272, 64'd3217477851037166, - 64'd3608713553388774, 64'd866972401106281, - 64'd146384793403658, 64'd6723655676905, 64'd152557945293083776, 64'd210512897111020, - 64'd3200744733577254, 64'd822260706595848, - 64'd149094118481168, 64'd9176796484705, 64'd151953595140331552, - 64'd2592926985077038, - 64'd2791379221130930, 64'd773084287120493, - 64'd150254851529169, 64'd11378404419023, 64'd150000908951494912, - 64'd5181109913618864, - 64'd2384456126063290, 64'd720197916448938, - 64'd149962184763602, 64'd13325531523291, 64'd146809868970192032, - 64'd7545074127449066, - 64'd1983529915919408, 64'd664338726404482, - 64'd148318097873735, 64'd15017758507562},
		'{64'd499867065461532032, - 64'd59090603245060688, 64'd13210686701393568, - 64'd2111808558266811, 64'd337486324545884, - 64'd46664229133003, 64'd470900528816664896, - 64'd56779642225398736, 64'd12665122499522302, - 64'd2055393536120170, 64'd331625184216959, - 64'd46986124451046, 64'd443082857930965312, - 64'd54496036558152024, 64'd12128490557472538, - 64'd1997406108287206, 64'd325205441481583, - 64'd47120469326447, 64'd416399082355731648, - 64'd52244856289559680, 64'd11601746744219710, - 64'd1938188289600451, 64'd318301134484187, - 64'd47084457892037, 64'd390831844704089728, - 64'd50030585969774272, 64'd11085723908655618, - 64'd1878054038124075, 64'd310980958127710, - 64'd46894236946073, 64'd366361683299355904, - 64'd47857164723061856, 64'd10581140665053968, - 64'd1817290843738338, 64'd303308536808829, - 64'd46564950434941, 64'd342967295276573248, - 64'd45728024374004640, 64'd10088609734400426, - 64'd1756161255870180, 64'd295342688467224, - 64'd46110783107821, 64'd320625781095457152, - 64'd43646125684975064, 64'd9608645855449780, - 64'd1694904350981282, 64'd287137679882200, - 64'd45545003275082, 64'd299312871395057152, - 64'd41613992761271952, 64'd9141673279508884, - 64'd1633737140569044, 64'd278743473185562, - 64'd44880004611618, 64'd279003137092026112, - 64'd39633745681138152, 64'd8688032863020428, - 64'd1572855920563987, 64'd270205963591973, - 64'd44127346955046, 64'd259670183595633024, - 64'd37707131408436864, 64'd8247988772044685, - 64'd1512437563120116, 64'd261567208377288, - 64'd43297796056757, 64'd241286829983672032, - 64'd35835553046077472, 64'd7821734812709202, - 64'd1452640751893828, 64'd252865647161803, - 64'd42401362251306, 64'd223825273954350464, - 64'd34020097488369872, 64'd7409400401624773, - 64'd1393607161993090, 64'd244136313579081, - 64'd41447338016438, 64'd207257243340165024, - 64'd32261561530372436, 64'd7011056190154086, - 64'd1335462585852560, 64'd235411038432292, - 64'd40444334402412, 64'd191554134940811712, - 64'd30560476492000676, 64'd6626719356271800, - 64'd1278318006353256, 64'd226718644458878, - 64'd39400316315058, 64'd176687141403401280, - 64'd28917131414200720, 64'd6256358577574866, - 64'd1222270618557855, 64'd218085132841096, - 64'd38322636642302, 64'd162627366849746080, - 64'd27331594883880184, 64'd5899898698793624, - 64'd1167404801475774, 64'd209533861614662, - 64'd37218069218740, 64'd149345931922318720, - 64'd25803735543545344, 64'd5557225106920785, - 64'd1113793041306316, 64'd201085716140550, - 64'd36092840627222, 64'd136814068892718880, - 64'd24333241340732608, 64'd5228187826820048, - 64'd1061496807634421, 64'd192759271815981, - 64'd34952660840432, 64'd125003207449179456, - 64'd22919637571358080, 64'd4912605349901751, - 64'd1010567384072244, 64'd184570949210115, - 64'd33802752709010, 64'd113885051752838192, - 64'd21562303770053916, 64'd4610268208162217, - 64'd961046654851821, 64'd176535161817829, - 64'd32647880306038, 64'd103431649326250800, - 64'd20260489499427320, 64'd4320942305578959, - 64'd912967848879905, 64'd168664456631467, - 64'd31492376140603, 64'd93615452311947264, - 64'd19013329088977392, 64'd4044372018537922, - 64'd866356242766271, 64'd160969647735727, - 64'd30340167255739, 64'd84409371613781216, - 64'd17819855373147846, 64'd3780283076643548, - 64'd821229824331948, 64'd153459943134852, - 64'd29194800228354, 64'd75786824409404512, - 64'd16679012476688924, 64'd3528385234929742, - 64'd777599918094377, 64'd146143065024310, - 64'd28059465090748},
		'{- 64'd499867065461795712, 64'd59090603245080680, - 64'd13210686701401844, 64'd2111808558268806, - 64'd337486324546168, 64'd46664229133005, - 64'd470900528816946240, 64'd56779642225419912, - 64'd12665122499531124, 64'd2055393536122300, - 64'd331625184217262, 64'd46986124451048, - 64'd443082857931261568, 64'd54496036558174208, - 64'd12128490557481822, 64'd1997406108289451, - 64'd325205441481902, 64'd47120469326449, - 64'd416399082356040512, 64'd52244856289582696, - 64'd11601746744229382, 64'd1938188289602794, - 64'd318301134484520, 64'd47084457892039, - 64'd390831844704409024, 64'd50030585969797968, - 64'd11085723908665608, 64'd1878054038126498, - 64'd310980958128054, 64'd46894236946075, - 64'd366361683299683520, 64'd47857164723086096, - 64'd10581140665064214, 64'd1817290843740825, - 64'd303308536809182, 64'd46564950434943, - 64'd342967295276907328, 64'd45728024374029288, - 64'd10088609734410870, 64'd1756161255872717, - 64'd295342688467585, 64'd46110783107823, - 64'd320625781095795968, 64'd43646125684999984, - 64'd9608645855460366, 64'd1694904350983856, - 64'd287137679882566, 64'd45545003275084, - 64'd299312871395399104, 64'd41613992761297056, - 64'd9141673279519566, 64'd1633737140571642, - 64'd278743473185931, 64'd44880004611621, - 64'd279003137092369760, 64'd39633745681163320, - 64'd8688032863031160, 64'd1572855920566600, - 64'd270205963592344, 64'd44127346955048, - 64'd259670183595977088, 64'd37707131408462016, - 64'd8247988772055426, 64'd1512437563122732, - 64'd261567208377660, 64'd43297796056759, - 64'd241286829984015296, 64'd35835553046102528, - 64'd7821734812719916, 64'd1452640751896438, - 64'd252865647162174, 64'd42401362251308, - 64'd223825273954691904, 64'd34020097488394756, - 64'd7409400401635427, 64'd1393607161995687, - 64'd244136313579450, 64'd41447338016440, - 64'd207257243340503616, 64'd32261561530397076, - 64'd7011056190164649, 64'd1335462585855137, - 64'd235411038432658, 64'd40444334402414, - 64'd191554134941146624, 64'd30560476492025016, - 64'd6626719356282246, 64'd1278318006355804, - 64'd226718644459240, 64'd39400316315060, - 64'd176687141403731680, 64'd28917131414224700, - 64'd6256358577585169, 64'd1222270618560370, - 64'd218085132841453, 64'd38322636642304, - 64'd162627366850071328, 64'd27331594883903768, - 64'd5899898698803765, 64'd1167404801478250, - 64'd209533861615014, 64'd37218069218742, - 64'd149345931922638208, 64'd25803735543568488, - 64'd5557225106930745, 64'd1113793041308748, - 64'd201085716140896, 64'd36092840627223, - 64'd136814068893032080, 64'd24333241340755272, - 64'd5228187826829810, 64'd1061496807636806, - 64'd192759271816320, 64'd34952660840433, - 64'd125003207449485904, 64'd22919637571380236, - 64'd4912605349911303, 64'd1010567384074578, - 64'd184570949210447, 64'd33802752709011, - 64'd113885051753137552, 64'd21562303770075536, - 64'd4610268208171545, 64'd961046654854101, - 64'd176535161818153, 64'd32647880306039, - 64'd103431649326542656, 64'd20260489499448380, - 64'd4320942305588053, 64'd912967848882128, - 64'd168664456631783, 64'd31492376140604, - 64'd93615452312231392, 64'd19013329088997876, - 64'd4044372018546774, 64'd866356242768436, - 64'd160969647736034, 64'd30340167255741, - 64'd84409371614057376, 64'd17819855373167740, - 64'd3780283076652152, 64'd821229824334052, - 64'd153459943135151, 64'd29194800228355, - 64'd75786824409672544, 64'd16679012476708220, - 64'd3528385234938091, 64'd777599918096419, - 64'd146143065024600, 64'd28059465090749}};
	localparam logic signed[63:0] Fbr[0:5][0:149] = '{
		'{64'd113364990210738416, - 64'd3983886949576016, - 64'd5569828753829607, - 64'd257905633687294, 64'd125531372261044, 64'd19081521365657, 64'd114421661700765920, - 64'd252787103572623, - 64'd5431958010978724, - 64'd364655848560909, 64'd112480991897162, 64'd20439689021416, 64'd113632587199134496, 64'd3389547035691944, - 64'd5211139927079489, - 64'd462952836698487, 64'd97966540628453, 64'd21439061241915, 64'd111056214328367104, 64'd6887404564960130, - 64'd4912948569680208, - 64'd551443750702659, 64'd82255227722555, 64'd22072669137832, 64'd106777957837526336, 64'd10188757390959440, - 64'd4544049735880285, - 64'd628965316574561, 64'd65626649275951, 64'd22339533300416, 64'd100908170763820064, 64'd13245995967219460, - 64'd4112067807347828, - 64'd694557617108024, 64'd48368034197952, 64'd22244530428458, 64'd93579769493015312, 64'd16016576473275068, - 64'd3625440673530840, - 64'd747474298852112, 64'd30769487045376, 64'd21798170151482, 64'd84945559090488032, 64'd18463571347437996, - 64'd3093265326712530, - 64'd787189129275752, 64'd13119303432000, 64'd21016287831245, 64'd75175308887683760, 64'd20556116822289656, - 64'd2525136816144404, - 64'd813398890629686, - 64'd4300569300313, 64'd19919660315895, 64'd64452631037034520, 64'd22269752907785916, - 64'd1930983287264629, - 64'd826022655588578, - 64'd21218857579341, 64'd18533552672876, 64'd52971716570588112, 64'd23586653090378920, - 64'd1320899826471287, - 64'd825197546169895, - 64'd37379009805054, 64'd16887204824597, 64'd40933984407312960, 64'd24495742838164032, - 64'd704983783260547, - 64'd811271130823059, - 64'd52542909780549, 64'd15013267744604, 64'd28544698759471100, 64'd24992707792833616, - 64'd93174151604766, - 64'd784790664188415, - 64'd66494204647644, 64'd12947199433882, 64'd16009609512006336, 64'd25079894261453868, 64'd504902536308573, - 64'd746489419146093, - 64'd79041203994704, 64'd10726631282315, 64'd3531668426439428, 64'd24766106268687644, 64'd1080077515416534, - 64'd697270400804040, - 64'd90019314700874, 64'd8390715627535, - 64'd8692128499272152, 64'd24066304968969788, 64'd1623774200497883, - 64'd638187766502393, - 64'd99292984344543, 64'd5979465353495, - 64'd20473725441161716, 64'd23001217626535588, 64'd2128129839791589, - 64'd570426304329795, - 64'd106757134494146, 64'd3533096228055, - 64'd31636774781455288, 64'd21596864629957068, 64'd2586102792344198, - 64'd495279344753834, - 64'd112338073775578, 64'd1091382369241, - 64'd42019150127781576, 64'd19884014100661044, 64'd2991564080733010, - 64'd414125495567832, - 64'd115993889134106, - 64'd1306965237301, - 64'd51475170700469208, 64'd17897574568536412, 64'd3339372154386992, - 64'd328404599363619, - 64'd117714322045471, - 64'd3624887860422, - 64'd59877508894710776, 64'd15675936912113984, 64'd3625430092182028, - 64'd239593315175250, - 64'd117520144452945, - 64'd5827527222024, - 64'd67118758563459712, 64'd13260277289108012, 64'd3846724771409130, - 64'd149180721926746, - 64'd115462056794691, - 64'd7882725072588, - 64'd73112647520344288, 64'd10693833111819658, 64'd4001347828734964, - 64'd58644331081793, - 64'd111619137529093, - 64'd9761467408887, - 64'd77794883829637216, 64'd8021164250755380, 64'd4088498532644028, 64'd30573120247393, - 64'd106096879966224, - 64'd11438267646808, - 64'd81123631533078432, 64'd5287411581728942, 64'd4108468971513664, 64'd117085746117695, - 64'd99024857885551, - 64'd12891484174376},
		'{64'd113364990210668768, - 64'd3983886949580926, - 64'd5569828753831866, - 64'd257905633687862, 64'd125531372260965, 64'd19081521365658, 64'd114421661700723616, - 64'd252787103575427, - 64'd5431958010980114, - 64'd364655848561268, 64'd112480991897113, 64'd20439689021417, 64'd113632587199119552, 64'd3389547035691238, - 64'd5211139927080010, - 64'd462952836698636, 64'd97966540628433, 64'd21439061241916, 64'd111056214328379040, 64'd6887404564961484, - 64'd4912948569679872, - 64'd551443750702600, 64'd82255227722564, 64'd22072669137833, 64'd106777957837564336, 64'd10188757390962776, - 64'd4544049735879120, - 64'd628965316574301, 64'd65626649275989, 64'd22339533300417, 64'd100908170763882864, 64'd13245995967224680, - 64'd4112067807345872, - 64'd694557617107572, 64'd48368034198017, 64'd22244530428459, 64'd93579769493101280, 64'd16016576473282042, - 64'd3625440673528145, - 64'd747474298851480, 64'd30769487045467, 64'd21798170151483, 64'd84945559090595232, 64'd18463571347446564, - 64'd3093265326709158, - 64'd787189129274954, 64'd13119303432114, 64'd21016287831246, 64'd75175308887809968, 64'd20556116822299648, - 64'd2525136816140422, - 64'd813398890628739, - 64'd4300569300178, 64'd19919660315896, 64'd64452631037177248, 64'd22269752907797136, - 64'd1930983287260118, - 64'd826022655587501, - 64'd21218857579189, 64'd18533552672878, 64'd52971716570744688, 64'd23586653090391160, - 64'd1320899826466332, - 64'd825197546168708, - 64'd37379009804886, 64'd16887204824598, 64'd40933984407480536, 64'd24495742838177072, - 64'd704983783255237, - 64'd811271130821784, - 64'd52542909780369, 64'd15013267744605, 64'd28544698759646752, 64'd24992707792847228, - 64'd93174151599195, - 64'd784790664187074, - 64'd66494204647454, 64'd12947199433883, 64'd16009609512187064, 64'd25079894261467816, 64'd504902536314311, - 64'd746489419144709, - 64'd79041203994508, 64'd10726631282316, 64'd3531668426622232, 64'd24766106268701704, 64'd1080077515422342, - 64'd697270400802637, - 64'd90019314700676, 64'd8390715627536, - 64'd8692128499090228, 64'd24066304968983732, 64'd1623774200503669, - 64'd638187766500992, - 64'd99292984344346, 64'd5979465353495, - 64'd20473725440983556, 64'd23001217626549200, 64'd2128129839797260, - 64'd570426304328420, - 64'd106757134493953, 64'd3533096228056, - 64'd31636774781283612, 64'd21596864629970132, 64'd2586102792349668, - 64'd495279344752505, - 64'd112338073775392, 64'd1091382369241, - 64'd42019150127618968, 64'd19884014100673372, 64'd2991564080738195, - 64'd414125495566571, - 64'd115993889133928, - 64'd1306965237301, - 64'd51475170700318016, 64'd17897574568547828, 64'd3339372154391818, - 64'd328404599362442, - 64'd117714322045306, - 64'd3624887860422, - 64'd59877508894573136, 64'd15675936912124328, 64'd3625430092186428, - 64'd239593315174175, - 64'd117520144452794, - 64'd5827527222024, - 64'd67118758563337464, 64'd13260277289117144, 64'd3846724771413042, - 64'd149180721925787, - 64'd115462056794557, - 64'd7882725072588, - 64'd73112647520238992, 64'd10693833111827464, 64'd4001347828738340, - 64'd58644331080962, - 64'd111619137528977, - 64'd9761467408887, - 64'd77794883829550112, 64'd8021164250761770, 64'd4088498532646828, 64'd30573120248085, - 64'd106096879966127, - 64'd11438267646808, - 64'd81123631533010496, 64'd5287411581733847, 64'd4108468971515856, 64'd117085746118241, - 64'd99024857885475, - 64'd12891484174376},
		'{64'd261185979523892064, - 64'd22456890558529396, - 64'd8607393505184881, - 64'd1769784954461006, - 64'd241447559502841, 64'd1933593015434, 64'd270800817222180096, - 64'd16047694531985916, - 64'd7900070649760353, - 64'd1716378903106676, - 64'd254857519535561, - 64'd3773288418972, 64'd277282227462791680, - 64'd9929647949627100, - 64'd7168828679240094, - 64'd1650925382366498, - 64'd265020553967774, - 64'd9055741381813, 64'd280785027968515808, - 64'd4138808128063452, - 64'd6421989129967633, - 64'd1574846110810426, - 64'd272065566502174, - 64'd13894456389570, 64'd281480698205836832, 64'd1294223557194100, - 64'd5667447612258315, - 64'd1489562841760350, - 64'd276141168090658, - 64'd18275501295111, 64'd279554672781074240, 64'd6344208747836490, - 64'd4912630705697034, - 64'd1396484358864565, - 64'd277412971381418, - 64'd22190081292982, 64'd275203692143743456, 64'd10991136482630424, - 64'd4164460088880028, - 64'd1296994478805553, - 64'd276060914540424, - 64'd25634268340864, 64'd268633230909669152, 64'd15220049038531744, - 64'd3429323737345382, - 64'd1192441102045094, - 64'd272276636914191, - 64'd28608704561309, 64'd260055022018696416, 64'd19020833458887984, - 64'd2713053970157080, - 64'd1084126340131656, - 64'd266260926991562, - 64'd31118284113950, 64'd249684692820901536, 64'd22387983019644088, - 64'd2020912077975607, - 64'd973297736300737, - 64'd258221261063288, - 64'd33171817918496, 64'd237739527061999296, 64'd25320332868942032, - 64'd1357579223514040, - 64'd861140584957512, - 64'd248369448891663, - 64'd34781685466361, 64'd224436364632737920, 64'd27820774022308884, - 64'd727153269036316, - 64'd748771345199828, - 64'd236919400609314, - 64'd35963477787308, 64'd209989648876552352, 64'd29895949807821008, - 64'd133151154946584, - 64'd637232133865376, - 64'd224085026986094, - 64'd36735635440535, 64'd194609629231121920, 64'd31555938736379624, 64'd421483571559838, - 64'd527486274706295, - 64'd210078283153949, - 64'd37119085180767, 64'd178500725027667200, 64'd32813927624776528, 64'd934368498510874, - 64'd420414872234720, - 64'd195107363878338, - 64'd37136878712585, 64'd161860054400109248, 64'd33685878626842608, 64'd1403665797068552, - 64'd316814371561296, - 64'd179375056526202, - 64'd36813836693955, 64'd144876130476242112, 64'd34190193633935372, 64'd1828061820100178, - 64'd217395059174395, - 64'd163077256018137, - 64'd36176200885914, 64'd127727725344849952, 64'd34347379293590144, 64'd2206743300987920, - 64'd122780454080956, - 64'd146401644278134, - 64'd35251297072942, 64'd110582900724628400, 64'd34179715667531056, 64'd2539370602628581, - 64'd33507534043250, - 64'd129526535018160, - 64'd34067211100752, 64'd93598202809657440, 64'd33710931310532892, 64'd2826048462808806, 64'd49972262215125, - 64'd112619883125651, - 64'd32652480097898, 64'd76918017437303328, 64'd32965887302861392, 64'd3067294674551256, 64'd127291319017218, - 64'd95838456466683, - 64'd31035800667583, 64'd60674080521596304, 64'd31970272514089748, 64'd3264007128945235, 64'd198163478416821, - 64'd79327166581764, - 64'd29245755558798, 64'd44985137620731944, 64'd30750312117747640, 64'd3417429633740691, 64'd262381091554607, - 64'd63218553538739, - 64'd27310560053785, 64'd29956745562421616, 64'd29332491117099896, 64'd3529116903943056, 64'd319811553507675, - 64'd47632419121166, - 64'd25257829044054, 64'd15681208235173768, 64'd27743294384802212, 64'd3600899101145688, 64'd370393388611762, - 64'd32675601571658, - 64'd23114365511491},
		'{64'd261185979523428576, - 64'd22456890558562344, - 64'd8607393505199444, - 64'd1769784954464604, - 64'd241447559503349, 64'd1933593015434, 64'd270800817221775808, - 64'd16047694532014440, - 64'd7900070649773052, - 64'd1716378903109822, - 64'd254857519536005, - 64'd3773288418972, 64'd277282227462446208, - 64'd9929647949651234, - 64'd7168828679250940, - 64'd1650925382369192, - 64'd265020553968155, - 64'd9055741381813, 64'd280785027968228288, - 64'd4138808128083280, - 64'd6421989129976653, - 64'd1574846110812677, - 64'd272065566502491, - 64'd13894456389570, 64'd281480698205605952, 64'd1294223557178464, - 64'd5667447612265551, - 64'd1489562841762165, - 64'd276141168090914, - 64'd18275501295111, 64'd279554672780898240, 64'd6344208747824902, - 64'd4912630705702542, - 64'd1396484358865959, - 64'd277412971381615, - 64'd22190081292981, 64'd275203692143620224, 64'd10991136482622716, - 64'd4164460088883876, - 64'd1296994478806542, - 64'd276060914540563, - 64'd25634268340863, 64'd268633230909596192, 64'd15220049038527722, - 64'd3429323737347648, - 64'd1192441102045696, - 64'd272276636914275, - 64'd28608704561307, 64'd260055022018670912, 64'd19020833458887424, - 64'd2713053970157851, - 64'd1084126340131892, - 64'd266260926991594, - 64'd31118284113949, 64'd249684692820920544, 64'd22387983019646772, - 64'd2020912077974979, - 64'd973297736300630, - 64'd258221261063272, - 64'd33171817918495, 64'd237739527062059552, 64'd25320332868947704, - 64'd1357579223512113, - 64'd861140584957086, - 64'd248369448891602, - 64'd34781685466359, 64'd224436364632836096, 64'd27820774022317292, - 64'd727153269033198, - 64'd748771345199110, - 64'd236919400609212, - 64'd35963477787306, 64'd209989648876684928, 64'd29895949807831892, - 64'd133151154942383, - 64'd637232133864391, - 64'd224085026985954, - 64'd36735635440533, 64'd194609629231285376, 64'd31555938736392708, 64'd421483571565008, - 64'd527486274705071, - 64'd210078283153775, - 64'd37119085180765, 64'd178500725027857888, 64'd32813927624791544, 64'd934368498516900, - 64'd420414872233284, - 64'd195107363878135, - 64'd37136878712583, 64'd161860054400323584, 64'd33685878626859292, 64'd1403665797075320, - 64'd316814371559676, - 64'd179375056525972, - 64'd36813836693953, 64'd144876130476476512, 64'd34190193633953452, 64'd1828061820107576, - 64'd217395059172618, - 64'd163077256017885, - 64'd36176200885912, 64'd127727725345100896, 64'd34347379293609364, 64'd2206743300995836, - 64'd122780454079049, - 64'd146401644277863, - 64'd35251297072941, 64'd110582900724892480, 64'd34179715667551152, 64'd2539370602636909, - 64'd33507534041241, - 64'd129526535017876, - 64'd34067211100751, 64'd93598202809931344, 64'd33710931310553636, 64'd2826048462817442, 64'd49972262217212, - 64'd112619883125355, - 64'd32652480097896, 64'd76918017437583840, 64'd32965887302882540, 64'd3067294674560098, 64'd127291319019360, - 64'd95838456466380, - 64'd31035800667582, 64'd60674080521880440, 64'd31970272514111080, 64'd3264007128954190, 64'd198163478418993, - 64'd79327166581456, - 64'd29245755558796, 64'd44985137621016856, 64'd30750312117768944, 64'd3417429633749668, 64'd262381091556787, - 64'd63218553538431, - 64'd27310560053784, 64'd29956745562704656, 64'd29332491117120984, 64'd3529116903951972, 64'd319811553509842, - 64'd47632419120859, - 64'd25257829044053, 64'd15681208235452464, 64'd27743294384822912, 64'd3600899101154465, 64'd370393388613898, - 64'd32675601571355, - 64'd23114365511490},
		'{64'd147927123522367456, - 64'd18177492446279264, - 64'd3137698184896970, - 64'd1488192028122724, - 64'd338884941609365, - 64'd83132750190217, 64'd156324607661916704, - 64'd15447556199019812, - 64'd2572490864587542, - 64'd1349781309511470, - 64'd311842990457516, - 64'd77626660430557, 64'd163408861711848480, - 64'd12922733796088518, - 64'd2051844969362986, - 64'd1219873695525226, - 64'd286301234270640, - 64'd72378730192471, 64'd169279715903773056, - 64'd10592180041143310, - 64'd1573311048560416, - 64'd1098104073152683, - 64'd262204033560234, - 64'd67382238575553, 64'd174031670337643904, - 64'd8445419759004248, - 64'd1134529129707866, - 64'd984114438549139, - 64'd239496148021515, - 64'd62630255352860, 64'd177754080110616032, - 64'd6472348047584440, - 64'd733228199975529, - 64'd877554426523398, - 64'd218122883876100, - 64'd58115683859598, 64'd180531340250850880, - 64'd4663229266772438, - 64'd367225438650931, - 64'd778081764645723, - 64'd198030225524146, - 64'd53831300404132, 64'd182443069855621344, - 64'd3008694886471708, - 64'd34425226629464, - 64'd685362657548161, - 64'd179164952541371, - 64'd49769790396593, 64'd183564294892240736, - 64'd1499740308324762, 64'd267182042787098, - 64'd599072106698097, - 64'd161474743008033, - 64'd45923781382925, 64'd183965629175753376, - 64'd127720768310654, 64'd539521329111766, - 64'd518894170645069, - 64'd144908264109849, - 64'd42285873164940, 64'd183713453089154848, 64'd1115653579602926, 64'd784434464784578, - 64'd444522170469735, - 64'd129415250904971, - 64'd38848665179692, 64'd182870089660314496, 64'd2238323305255050, 64'd1003681810516536, - 64'd375658844902448, - 64'd114946574106669, - 64'd35604781304352, 64'd181493977654918944, 64'd3247885982404254, 64'd1198944027602716, - 64'd312016459327057, - 64'd101454297688191, - 64'd32546892245770, 64'd179639841386790816, 64'd4151603026088577, 64'd1371823950268495, - 64'd253316872643342, - 64'd88891727074462, - 64'd29667735666990, 64'd177358856986020544, 64'd4956407011924468, 64'd1523848542371368, - 64'd199291565728716, - 64'd77213448644859, - 64'd26960134196258, 64'd174698814901622912, 64'd5668909407507587, 64'd1656470923973247, - 64'd149681635016508, - 64'd66375361232269, - 64'd24417011457433, 64'd171704278449040032, 64'd6295408651269154, 64'd1771072454427026, - 64'd104237754493935, - 64'd56334700265924, - 64'd22031406254313, 64'd168416738243893632, 64'd6841898519060024, 64'd1868964859688488, - 64'd62720109217924, - 64'd47050055169258, - 64'd19796485035030, 64'd164874762392079616, 64'd7314076723390628, 64'd1951392392572694, - 64'd24898303250727, - 64'd38481380589084, - 64'd17705552756628, 64'd161114142332723552, 64'd7717353694656953, 64'd2019534015624960, 64'd9448755270026, - 64'd30590001998816, - 64'd15752062263952, 64'd157168034254798720, 64'd8056861497840441, 64'd2074505597172628, 64'd40532989391103, - 64'd23338616186249, - 64'd13929622291208, 64'd153067096030477760, 64'd8337462842091858, 64'd2117362111967220, 64'd68557306567997, - 64'd16691287105506, - 64'd12232004189014, 64'd148839619628647360, 64'd8563760144304924, 64'd2149099838619291, 64'd93715767650942, - 64'd10613437543130, - 64'd10653147474290, 64'd144511658990586496, 64'd8740104611263724, 64'd2170658546772659, 64'd116193769584212, - 64'd5071837020033, - 64'd9187164295181, 64'd140107153366689824, 64'd8870605308217606, 64'd2182923667662533, 64'd136168239917123, - 64'd34586323870, - 64'd7828342898123},
		'{64'd147927123521392000, - 64'd18177492446348480, - 64'd3137698184927293, - 64'd1488192028130171, - 64'd338884941610422, - 64'd83132750190221, 64'd156324607660996992, - 64'd15447556199085032, - 64'd2572490864616129, - 64'd1349781309518492, - 64'd311842990458513, - 64'd77626660430561, 64'd163408861710982336, - 64'd12922733796149900, - 64'd2051844969389905, - 64'd1219873695531840, - 64'd286301234271579, - 64'd72378730192475, 64'd169279715902958368, - 64'd10592180041201008, - 64'd1573311048585734, - 64'd1098104073158904, - 64'd262204033561118, - 64'd67382238575556, 64'd174031670336878528, - 64'd8445419759058417, - 64'd1134529129731650, - 64'd984114438554984, - 64'd239496148022345, - 64'd62630255352863, 64'd177754080109897920, - 64'd6472348047635232, - 64'd733228199997842, - 64'd877554426528883, - 64'd218122883876879, - 64'd58115683859601, 64'd180531340250177952, - 64'd4663229266820000, - 64'd367225438671837, - 64'd778081764650863, - 64'd198030225524876, - 64'd53831300404135, 64'd182443069854991616, - 64'd3008694886516184, - 64'd34425226649026, - 64'd685362657552972, - 64'd179164952542054, - 64'd49769790396595, 64'd183564294891652288, - 64'd1499740308366294, 64'd267182042768819, - 64'd599072106702593, - 64'd161474743008671, - 64'd45923781382927, 64'd183965629175204256, - 64'd127720768349380, 64'd539521329094712, - 64'd518894170649265, - 64'd144908264110445, - 64'd42285873164942, 64'd183713453088643200, 64'd1115653579566872, 64'd784434464768689, - 64'd444522170473645, - 64'd129415250905526, - 64'd38848665179694, 64'd182870089659838528, 64'd2238323305221536, 64'd1003681810501757, - 64'd375658844906086, - 64'd114946574107185, - 64'd35604781304353, 64'd181493977654476864, 64'd3247885982373158, 64'd1198944027588991, - 64'd312016459330436, - 64'd101454297688671, - 64'd32546892245771, 64'd179639841386380928, 64'd4151603026059772, 64'd1371823950255771, - 64'd253316872646475, - 64'd88891727074907, - 64'd29667735666992, 64'd177358856985641184, 64'd4956407011897833, 64'd1523848542359593, - 64'd199291565731617, - 64'd77213448645271, - 64'd26960134196259, 64'd174698814901272480, 64'd5668909407483011, 64'd1656470923962372, - 64'd149681635019187, - 64'd66375361232649, - 64'd24417011457435, 64'd171704278448716992, 64'd6295408651246523, 64'd1771072454417002, - 64'd104237754496406, - 64'd56334700266274, - 64'd22031406254314, 64'd168416738243596480, 64'd6841898519039232, 64'd1868964859679269, - 64'd62720109220197, - 64'd47050055169581, - 64'd19796485035031, 64'd164874762391806912, 64'd7314076723371573, 64'd1951392392564236, - 64'd24898303252813, - 64'd38481380589380, - 64'd17705552756629, 64'd161114142332473920, 64'd7717353694639534, 64'd2019534015617218, 64'd9448755268116, - 64'd30590001999087, - 64'd15752062263952, 64'd157168034254570816, 64'd8056861497824561, 64'd2074505597165561, 64'd40532989389359, - 64'd23338616186497, - 64'd13929622291209, 64'd153067096030270272, 64'd8337462842077426, 64'd2117362111960788, 64'd68557306566409, - 64'd16691287105731, - 64'd12232004189015, 64'd148839619628459104, 64'd8563760144291853, 64'd2149099838613457, 64'd93715767649500, - 64'd10613437543335, - 64'd10653147474290, 64'd144511658990416288, 64'd8740104611251929, 64'd2170658546767385, 64'd116193769582909, - 64'd5071837020218, - 64'd9187164295182, 64'd140107153366536528, 64'd8870605308207004, 64'd2182923667657784, 64'd136168239915949, - 64'd34586324037, - 64'd7828342898124}};
	localparam logic signed[63:0] Fbi[0:5][0:149] = '{
		'{- 64'd27061454864742516, - 64'd29329963185269764, - 64'd195520791088329, 64'd900075992202870, 64'd84307738655099, - 64'd14039756020202, - 64'd12402408768204324, - 64'd29227842841782012, - 64'd884657663660782, 64'd849633769750120, 64'd98210562395013, - 64'd11379009668686, 64'd2089310716763816, - 64'd28663497405476736, - 64'd1542589681822757, 64'd786935553955462, 64'd110205960410614, - 64'd8603488459578, 64'd16187425555932316, - 64'd27657395440758048, - 64'd2159630788206751, 64'd713283119733266, 64'd120150622728524, - 64'd5760181395202, 64'd29677543699628088, - 64'd26236521060170792, - 64'd2726986023501624, 64'd630120057110324, 64'd127937412862532, - 64'd2895986842769, 64'd42360272641980240, - 64'd24433782808960836, - 64'd3236869219002734, 64'd539005289400233, 64'd133496171871328, - 64'd56969036973, 64'd54054017037580968, - 64'd22287343042577064, - 64'd3682601721153442, 64'd441585415965900, 64'd136793914424840, 64'd2712353664127, 64'd64597423746336640, - 64'd19839880438164920, - 64'd4058691049914580, 64'd339566348590174, 64'd137834428881022, 64'd5369678241846, 64'd73851444194581232, - 64'd17137799030007612, - 64'd4360888739188662, 64'd234684710043639, 64'd136657302553573, 64'd7875534604264, 64'd81700990774571280, - 64'd14230397676234388, - 64'd4586226957255934, 64'd128679455567068, 64'd133336401964652, 64'd10193842767793, 64'd88056171038730048, - 64'd11169014147466116, - 64'd4733033852605743, 64'd23264162984228, 64'd127977845802236, 64'd12292402275104, 64'd92853090562627088, - 64'd8006158078720994, - 64'd4800927910201560, - 64'd79899584555584, 64'd120717515430476, 64'd14143307752129, 64'd96054222436410784, - 64'd4794646848838514, - 64'd4790791929893918, - 64'd179227327124325, 64'd111718154039706, 64'd15723285832956, 64'd97648348286379680, - 64'd1586758055376818, - 64'd4704727547520385, - 64'd273235005292775, 64'd101166110793507, 64'd17013950050470, 64'd97650082419767936, 64'd1566588350849615, - 64'd4545991505738860, - 64'd360560062034348, 64'd89267790573839, 64'd18001971679645, 64'd96098997026461056, 64'd4616606003936770, - 64'd4318915141828897, - 64'd439980087802016, 64'd76245873099580, 64'd18679165906927, 64'd93058372269148240, 64'd7517364837884810, - 64'd4028808790082756, - 64'd510428773391513, 64'd62335367275175, 64'd19042494061181, 64'd88613600465584832, 64'd10226450409772886, - 64'd3681852994070874, - 64'd571008983867665, 64'd47779567608419, 64'd19093983958108, 64'd82870278340830400, 64'd12705550923365190, - 64'd3284978586676226, - 64'd621002817253347, 64'd32825979431485, 64'd18840571661139, 64'd75952025442497056, 64'd14920964416583992, - 64'd2845737821634594, - 64'd659878563016750, 64'd17722278495844, 64'd18293869129252, 64'd67998070219142936, 64'd16844020033214614, - 64'd2372168828306202, - 64'd687294526803150, 64'd2712368334485, 64'd17469863289503, 64'd59160647924404656, 64'd18451408816580252, - 64'd1872655711080900, - 64'd703099738523027, - 64'd11967404346242, 64'd16388553024781, 64'd49602256403463392, 64'd19725421015109816, - 64'd1355786626346778, - 64'd707331610041940, - 64'd26091819994366, 64'd15073531393143, 64'd39492816932973920, 64'd20654088451171928, - 64'd830212144096177, - 64'd700210655575872, - 64'd39450090815028, 64'd13551521084012, 64'd29006787622315340, 64'd21231232050203092, - 64'd304506139344359, - 64'd682132431790285, - 64'd51848853708365, 64'd11851871661078},
		'{64'd27061454864950924, 64'd29329963185285884, 64'd195520791094942, - 64'd900075992201277, - 64'd84307738654874, 64'd14039756020203, 64'd12402408768417152, 64'd29227842841798412, 64'd884657663667541, - 64'd849633769748489, - 64'd98210562394782, 64'd11379009668687, - 64'd2089310716550064, 64'd28663497405493156, 64'd1542589681829552, - 64'd786935553953819, - 64'd110205960410382, 64'd8603488459578, - 64'd16187425555721056, 64'd27657395440774216, 64'd2159630788213471, - 64'd713283119731638, - 64'd120150622728295, 64'd5760181395203, - 64'd29677543699422628, 64'd26236521060186464, 64'd2726986023508166, - 64'd630120057108737, - 64'd127937412862309, 64'd2895986842770, - 64'd42360272641783696, 64'd24433782808975776, 64'd3236869219008998, - 64'd539005289398711, - 64'd133496171871114, 64'd56969036974, - 64'd54054017037396248, 64'd22287343042591052, 64'd3682601721159334, - 64'd441585415964465, - 64'd136793914424639, - 64'd2712353664127, - 64'd64597423746166368, 64'd19839880438177752, 64'd4058691049920017, - 64'd339566348588847, - 64'd137834428880836, - 64'd5369678241846, - 64'd73851444194427808, 64'd17137799030019116, 64'd4360888739193568, - 64'd234684710042438, - 64'd136657302553405, - 64'd7875534604264, - 64'd81700990774436672, 64'd14230397676244412, 64'd4586226957260245, - 64'd128679455566009, - 64'd133336401964504, - 64'd10193842767793, - 64'd88056171038615952, 64'd11169014147474542, 64'd4733033852609405, - 64'd23264162983325, - 64'd127977845802110, - 64'd12292402275104, - 64'd92853090562534800, 64'd8006158078727724, 64'd4800927910204531, 64'd79899584556320, - 64'd120717515430374, - 64'd14143307752129, - 64'd96054222436341232, 64'd4794646848843485, 64'd4790791929896167, 64'd179227327124888, - 64'd111718154039628, - 64'd15723285832956, - 64'd97648348286333408, 64'd1586758055379994, 64'd4704727547521895, 64'd273235005293160, - 64'd101166110793454, - 64'd17013950050471, - 64'd97650082419745088, - 64'd1566588350848240, 64'd4545991505739625, 64'd360560062034553, - 64'd89267790573811, - 64'd18001971679646, - 64'd96098997026461440, - 64'd4616606003937172, 64'd4318915141828924, 64'd439980087802041, - 64'd76245873099577, - 64'd18679165906928, - 64'd93058372269171232, - 64'd7517364837886940, 64'd4028808790082064, 64'd510428773391364, - 64'd62335367275197, - 64'd19042494061182, - 64'd88613600465629536, - 64'd10226450409776666, 64'd3681852994069489, 64'd571008983867348, - 64'd47779567608464, - 64'd19093983958110, - 64'd82870278340895552, - 64'd12705550923370520, 64'd3284978586674188, 64'd621002817252871, - 64'd32825979431553, - 64'd18840571661141, - 64'd75952025442581120, - 64'd14920964416590748, 64'd2845737821631954, 64'd659878563016127, - 64'd17722278495933, - 64'd18293869129253, - 64'd67998070219244096, - 64'd16844020033222652, 64'd2372168828303015, 64'd687294526802393, - 64'd2712368334593, - 64'd17469863289504, - 64'd59160647924520880, - 64'd18451408816589412, 64'd1872655711077230, 64'd703099738522152, 64'd11967404346118, - 64'd16388553024782, - 64'd49602256403592464, - 64'd19725421015119928, 64'd1355786626342696, 64'd707331610040964, 64'd26091819994228, - 64'd15073531393144, - 64'd39492816933113472, - 64'd20654088451182804, 64'd830212144091758, 64'd700210655574812, 64'd39450090814878, - 64'd13551521084013, - 64'd29006787622462876, - 64'd21231232050214544, 64'd304506139339682, 64'd682132431789160, 64'd51848853708206, - 64'd11851871661079},
		'{- 64'd225677438598042560, - 64'd63354485394154200, - 64'd4276556762928860, 64'd173233147734769, 64'd260338546982839, 64'd64414188308395, - 64'd194099328777530528, - 64'd62863947226030400, - 64'd4863482625348990, 64'd11783768817828, 64'd229143648540106, 64'd62088170629478, - 64'd162903732143129920, - 64'd61832029002577360, - 64'd5365829956533783, - 64'd138742379771980, 64'd197984597261583, 64'd59353276176248, - 64'd132349799862027520, - 64'd60305157375926432, - 64'd5784783558645604, - 64'd277715051368705, 64'd167143895985067, 64'd56262452200578, - 64'd102673108580712048, - 64'd58331113296847152, - 64'd6122209925009098, - 64'd404652718271066, 64'd136881834266162, 64'd52868283349588, - 64'd74085116781183136, - 64'd55958502521860016, - 64'd6380593594475096, - 64'd519216814161826, 64'd107435625726572, 64'd49222535549607, - 64'd46772878844103376, - 64'd53236254754919808, - 64'd6562972202281639, - 64'd621205062519008, 64'd79018815374206, 64'd45375738541443, - 64'd20899001826037872, - 64'd50213154047608856, - 64'd6672870910438875, - 64'd710544014480569, 64'd51820943869420, 64'd41376808243854, 64'd3398171237329920, - 64'd46937402616638520, - 64'd6714236859671300, - 64'd787280918418317, 64'd26007454251939, 64'd37272709677485, 64'd26004168655667776, - 64'd43456219784353120, - 64'd6691374240886772, - 64'd851575041235286, 64'd1719825415355, 64'd33108160760582, 64'd46827805932517792, - 64'd39815477310187040, - 64'd6608880537620060, - 64'd903688558214912, - 64'd20924084383897, 64'd28925376892742, 64'd65800428562538304, - 64'd36059371961594712, - 64'd6471584442512415, - 64'd943977124213681, - 64'd41829501475068, 64'd24763855875645, 64'd82875000525838496, - 64'd32230135774440352, - 64'd6284485901207953, - 64'd972880234196613, - 64'd60924026236796, 64'd20660202381705, 64'd98025057357911808, - 64'd28367784077415996, - 64'd6052698686615020, - 64'd990911475662388, - 64'd78156766495518, 64'd16647990873758, 64'd111243542622272928, - 64'd24509901004605992, - 64'd5781395855809029, - 64'd998648769487086, - 64'd93497333446865, 64'd12757665602248, 64'd122541546392837312, - 64'd20691461896333824, - 64'd5475758391422012, - 64'd996724689226150, - 64'd106934718675527, 64'd9016476061142, 64'd131946963977888080, - 64'd16944691692066244, - 64'd5140927279618252, - 64'd985816942044687, - 64'd118476070667219, 64'd5448446070101, 64'd139503092601186624, - 64'd13298958151233642, - 64'd4781959228102836, - 64'd966639087285579, - 64'd128145388868866, 64'd2074374468180, 64'd145267183112758496, - 64'd9780698498861298, - 64'd4403786180421141, - 64'd939931561318297, - 64'd135982152873408, - 64'd1088134747168, 64'd149308963046665856, - 64'd6413377883100207, - 64'd4011178737413532, - 64'd906453069820362, - 64'd142039903698047, - 64'd4024615123238, 64'd151709146490235968, - 64'd3217477851025686, - 64'd3608713553383575, - 64'd866972401104986, - 64'd146384793403475, - 64'd6723655676905, 64'd152557945293218496, - 64'd210512897101834, - 64'd3200744733573030, - 64'd822260706594790, - 64'd149094118481018, - 64'd9176796484705, 64'd151953595140436224, 64'd2592926985084004, - 64'd2791379221127652, - 64'd773084287119666, - 64'd150254851529052, - 64'd11378404419024, 64'd150000908951570592, 64'd5181109913623697, - 64'd2384456126060925, - 64'd720197916448334, - 64'd149962184763518, - 64'd13325531523291, 64'd146809868970240064, 64'd7545074127451866, - 64'd1983529915917913, - 64'd664338726404090, - 64'd148318097873680, - 64'd15017758507562},
		'{64'd225677438598514048, 64'd63354485394190232, 64'd4276556762943734, - 64'd173233147731185, - 64'd260338546982331, - 64'd64414188308392, 64'd194099328778024256, 64'd62863947226067920, 64'd4863482625364560, - 64'd11783768814068, - 64'd229143648539574, - 64'd62088170629475, 64'd162903732143639872, 64'd61832029002615920, 64'd5365829956549861, 64'd138742379775869, - 64'd197984597261032, - 64'd59353276176245, 64'd132349799862547968, 64'd60305157375965608, 64'd5784783558662007, 64'd277715051372679, - 64'd167143895984504, - 64'd56262452200575, 64'd102673108581237456, 64'd58331113296886536, 64'd6122209925025654, 64'd404652718275083, - 64'd136881834265593, - 64'd52868283349585, 64'd74085116781708352, 64'd55958502521899248, 64'd6380593594491644, 64'd519216814165847, - 64'd107435625726003, - 64'd49222535549604, 64'd46772878844623648, 64'd53236254754958536, 64'd6562972202298028, 64'd621205062522994, - 64'd79018815373642, - 64'd45375738541441, 64'd20899001826548768, 64'd50213154047646760, 64'd6672870910454965, 64'd710544014484487, - 64'd51820943868866, - 64'd41376808243852, - 64'd3398171236832432, 64'd46937402616675296, 64'd6714236859686965, 64'd787280918422136, - 64'd26007454251399, - 64'd37272709677482, - 64'd26004168655187328, 64'd43456219784388528, 64'd6691374240901898, 64'd851575041238978, - 64'd1719825414833, - 64'd33108160760581, - 64'd46827805932057600, 64'd39815477310220848, 64'd6608880537634544, 64'd903688558218452, 64'd20924084384398, - 64'd28925376892740, - 64'd65800428562101232, 64'd36059371961626704, 64'd6471584442526171, 64'd943977124217046, 64'd41829501475544, - 64'd24763855875643, - 64'd82875000525426944, 64'd32230135774470372, 64'd6284485901220903, 64'd972880234199785, 64'd60924026237245, - 64'd20660202381703, - 64'd98025057357527776, 64'd28367784077443900, 64'd6052698686627101, 64'd990911475665351, 64'd78156766495936, - 64'd16647990873756, - 64'd111243542621918048, 64'd24509901004631672, 64'd5781395855820190, 64'd998648769489827, 64'd93497333447253, - 64'd12757665602247, - 64'd122541546392512864, 64'd20691461896357200, 64'd5475758391432213, 64'd996724689228659, 64'd106934718675882, - 64'd9016476061141, - 64'd131946963977594928, 64'd16944691692087254, 64'd5140927279627466, 64'd985816942046958, 64'd118476070667540, - 64'd5448446070100, - 64'd139503092600925328, 64'd13298958151252256, 64'd4781959228111047, 64'd966639087287606, 64'd128145388869152, - 64'd2074374468179, - 64'd145267183112529280, 64'd9780698498877512, 64'd4403786180428342, 64'd939931561320079, 64'd135982152873659, 64'd1088134747169, - 64'd149308963046468608, 64'd6413377883114036, 64'd4011178737419725, 64'd906453069821900, 64'd142039903698264, 64'd4024615123238, - 64'd151709146490070272, 64'd3217477851037166, 64'd3608713553388774, 64'd866972401106281, 64'd146384793403658, 64'd6723655676905, - 64'd152557945293083776, 64'd210512897111020, 64'd3200744733577254, 64'd822260706595848, 64'd149094118481168, 64'd9176796484705, - 64'd151953595140331552, - 64'd2592926985077038, 64'd2791379221130930, 64'd773084287120493, 64'd150254851529169, 64'd11378404419023, - 64'd150000908951494912, - 64'd5181109913618864, 64'd2384456126063290, 64'd720197916448938, 64'd149962184763602, 64'd13325531523291, - 64'd146809868970192032, - 64'd7545074127449066, 64'd1983529915919408, 64'd664338726404482, 64'd148318097873735, 64'd15017758507562},
		'{- 64'd499867065461532032, - 64'd59090603245060688, - 64'd13210686701393568, - 64'd2111808558266811, - 64'd337486324545884, - 64'd46664229133003, - 64'd470900528816664896, - 64'd56779642225398736, - 64'd12665122499522302, - 64'd2055393536120170, - 64'd331625184216959, - 64'd46986124451046, - 64'd443082857930965312, - 64'd54496036558152024, - 64'd12128490557472538, - 64'd1997406108287206, - 64'd325205441481583, - 64'd47120469326447, - 64'd416399082355731648, - 64'd52244856289559680, - 64'd11601746744219710, - 64'd1938188289600451, - 64'd318301134484187, - 64'd47084457892037, - 64'd390831844704089728, - 64'd50030585969774272, - 64'd11085723908655618, - 64'd1878054038124075, - 64'd310980958127710, - 64'd46894236946073, - 64'd366361683299355904, - 64'd47857164723061856, - 64'd10581140665053968, - 64'd1817290843738338, - 64'd303308536808829, - 64'd46564950434941, - 64'd342967295276573248, - 64'd45728024374004640, - 64'd10088609734400426, - 64'd1756161255870180, - 64'd295342688467224, - 64'd46110783107821, - 64'd320625781095457152, - 64'd43646125684975064, - 64'd9608645855449780, - 64'd1694904350981282, - 64'd287137679882200, - 64'd45545003275082, - 64'd299312871395057152, - 64'd41613992761271952, - 64'd9141673279508884, - 64'd1633737140569044, - 64'd278743473185562, - 64'd44880004611618, - 64'd279003137092026112, - 64'd39633745681138152, - 64'd8688032863020428, - 64'd1572855920563987, - 64'd270205963591973, - 64'd44127346955046, - 64'd259670183595633024, - 64'd37707131408436864, - 64'd8247988772044685, - 64'd1512437563120116, - 64'd261567208377288, - 64'd43297796056757, - 64'd241286829983672032, - 64'd35835553046077472, - 64'd7821734812709202, - 64'd1452640751893828, - 64'd252865647161803, - 64'd42401362251306, - 64'd223825273954350464, - 64'd34020097488369872, - 64'd7409400401624773, - 64'd1393607161993090, - 64'd244136313579081, - 64'd41447338016438, - 64'd207257243340165024, - 64'd32261561530372436, - 64'd7011056190154086, - 64'd1335462585852560, - 64'd235411038432292, - 64'd40444334402412, - 64'd191554134940811712, - 64'd30560476492000676, - 64'd6626719356271800, - 64'd1278318006353256, - 64'd226718644458878, - 64'd39400316315058, - 64'd176687141403401280, - 64'd28917131414200720, - 64'd6256358577574866, - 64'd1222270618557855, - 64'd218085132841096, - 64'd38322636642302, - 64'd162627366849746080, - 64'd27331594883880184, - 64'd5899898698793624, - 64'd1167404801475774, - 64'd209533861614662, - 64'd37218069218740, - 64'd149345931922318720, - 64'd25803735543545344, - 64'd5557225106920785, - 64'd1113793041306316, - 64'd201085716140550, - 64'd36092840627222, - 64'd136814068892718880, - 64'd24333241340732608, - 64'd5228187826820048, - 64'd1061496807634421, - 64'd192759271815981, - 64'd34952660840432, - 64'd125003207449179456, - 64'd22919637571358080, - 64'd4912605349901751, - 64'd1010567384072244, - 64'd184570949210115, - 64'd33802752709010, - 64'd113885051752838192, - 64'd21562303770053916, - 64'd4610268208162217, - 64'd961046654851821, - 64'd176535161817829, - 64'd32647880306038, - 64'd103431649326250800, - 64'd20260489499427320, - 64'd4320942305578959, - 64'd912967848879905, - 64'd168664456631467, - 64'd31492376140603, - 64'd93615452311947264, - 64'd19013329088977392, - 64'd4044372018537922, - 64'd866356242766271, - 64'd160969647735727, - 64'd30340167255739, - 64'd84409371613781216, - 64'd17819855373147846, - 64'd3780283076643548, - 64'd821229824331948, - 64'd153459943134852, - 64'd29194800228354, - 64'd75786824409404512, - 64'd16679012476688924, - 64'd3528385234929742, - 64'd777599918094377, - 64'd146143065024310, - 64'd28059465090748},
		'{64'd499867065461795712, 64'd59090603245080680, 64'd13210686701401844, 64'd2111808558268806, 64'd337486324546168, 64'd46664229133005, 64'd470900528816946240, 64'd56779642225419912, 64'd12665122499531124, 64'd2055393536122300, 64'd331625184217262, 64'd46986124451048, 64'd443082857931261568, 64'd54496036558174208, 64'd12128490557481822, 64'd1997406108289451, 64'd325205441481902, 64'd47120469326449, 64'd416399082356040512, 64'd52244856289582696, 64'd11601746744229382, 64'd1938188289602794, 64'd318301134484520, 64'd47084457892039, 64'd390831844704409024, 64'd50030585969797968, 64'd11085723908665608, 64'd1878054038126498, 64'd310980958128054, 64'd46894236946075, 64'd366361683299683520, 64'd47857164723086096, 64'd10581140665064214, 64'd1817290843740825, 64'd303308536809182, 64'd46564950434943, 64'd342967295276907328, 64'd45728024374029288, 64'd10088609734410870, 64'd1756161255872717, 64'd295342688467585, 64'd46110783107823, 64'd320625781095795968, 64'd43646125684999984, 64'd9608645855460366, 64'd1694904350983856, 64'd287137679882566, 64'd45545003275084, 64'd299312871395399104, 64'd41613992761297056, 64'd9141673279519566, 64'd1633737140571642, 64'd278743473185931, 64'd44880004611621, 64'd279003137092369760, 64'd39633745681163320, 64'd8688032863031160, 64'd1572855920566600, 64'd270205963592344, 64'd44127346955048, 64'd259670183595977088, 64'd37707131408462016, 64'd8247988772055426, 64'd1512437563122732, 64'd261567208377660, 64'd43297796056759, 64'd241286829984015296, 64'd35835553046102528, 64'd7821734812719916, 64'd1452640751896438, 64'd252865647162174, 64'd42401362251308, 64'd223825273954691904, 64'd34020097488394756, 64'd7409400401635427, 64'd1393607161995687, 64'd244136313579450, 64'd41447338016440, 64'd207257243340503616, 64'd32261561530397076, 64'd7011056190164649, 64'd1335462585855137, 64'd235411038432658, 64'd40444334402414, 64'd191554134941146624, 64'd30560476492025016, 64'd6626719356282246, 64'd1278318006355804, 64'd226718644459240, 64'd39400316315060, 64'd176687141403731680, 64'd28917131414224700, 64'd6256358577585169, 64'd1222270618560370, 64'd218085132841453, 64'd38322636642304, 64'd162627366850071328, 64'd27331594883903768, 64'd5899898698803765, 64'd1167404801478250, 64'd209533861615014, 64'd37218069218742, 64'd149345931922638208, 64'd25803735543568488, 64'd5557225106930745, 64'd1113793041308748, 64'd201085716140896, 64'd36092840627223, 64'd136814068893032080, 64'd24333241340755272, 64'd5228187826829810, 64'd1061496807636806, 64'd192759271816320, 64'd34952660840433, 64'd125003207449485904, 64'd22919637571380236, 64'd4912605349911303, 64'd1010567384074578, 64'd184570949210447, 64'd33802752709011, 64'd113885051753137552, 64'd21562303770075536, 64'd4610268208171545, 64'd961046654854101, 64'd176535161818153, 64'd32647880306039, 64'd103431649326542656, 64'd20260489499448380, 64'd4320942305588053, 64'd912967848882128, 64'd168664456631783, 64'd31492376140604, 64'd93615452312231392, 64'd19013329088997876, 64'd4044372018546774, 64'd866356242768436, 64'd160969647736034, 64'd30340167255741, 64'd84409371614057376, 64'd17819855373167740, 64'd3780283076652152, 64'd821229824334052, 64'd153459943135151, 64'd29194800228355, 64'd75786824409672544, 64'd16679012476708220, 64'd3528385234938091, 64'd777599918096419, 64'd146143065024600, 64'd28059465090749}};
	localparam logic signed[63:0] hf[0:1799] = {64'd11671469817856, - 64'd68906754048, - 64'd75389681664, 64'd632993600, 64'd1232912256, - 64'd13692950, 64'd11602687426560, - 64'd205972455424, - 64'd73580404736, 64'd1884879744, 64'd1207679872, - 64'd40773932, 64'd11465870278656, - 64'd340804698112, - 64'd69988712448, 64'd3094723328, 64'd1157783296, - 64'd66948644, 64'd11262497914880, - 64'd471947444224, - 64'd64667860992, 64'd4235354880, 64'd1084343936, - 64'd91640440, 64'd10994772344832, - 64'd597993521152, - 64'd57696690176, 64'd5280870912, 64'd989008640, - 64'd114312056, 64'd10665578201088, - 64'd717603078144, - 64'd49178345472, 64'd6207100416, 64'd873910592, - 64'd134478512, 64'd10278451281920, - 64'd829521199104, - 64'd39238668288, 64'd6992039424, 64'd741620736, - 64'd151718128, 64'd9837531365376, - 64'd932594057216, - 64'd28024207360, 64'd7616239104, 64'd595090240, - 64'd165681392, 64'd9347505586176, - 64'd1025783496704, - 64'd15699915776, 64'd8063150592, 64'd437586208, - 64'd176098000, 64'd8813547618304, - 64'd1108180467712, - 64'd2446590720, 64'd8319411200, 64'd272621824, - 64'd182781520, 64'd8241252663296, - 64'd1179015708672, 64'd11541940224, 64'd8375070720, 64'd103882200, - 64'd185632240, 64'd7636563001344, - 64'd1237668986880, 64'd26061805568, 64'd8223759872, - 64'd64851640, - 64'd184637792, 64'd7005691969536, - 64'd1283676045312, 64'd40902221824, 64'd7862790656, - 64'd229779984, - 64'd179871936, 64'd6355046367232, - 64'd1316733190144, 64'd55848693760, 64'd7293190144, - 64'd387160704, - 64'd171491536, 64'd5691141521408, - 64'd1336699518976, 64'd70686261248, 64'd6519671296, - 64'd533383328, - 64'd159731776, 64'd5020525789184, - 64'd1343597314048, 64'd85202714624, 64'd5550539264, - 64'd665039680, - 64'd144899840, 64'd4349692739584, - 64'd1337609420800, 64'd99191758848, 64'd4397536256, - 64'd778989504, - 64'd127367376, 64'd3685008015360, - 64'd1319074791424, 64'd112455999488, 64'd3075626240, - 64'd872420032, - 64'd107561680, 64'd3032628592640, - 64'd1288481931264, 64'd124809854976, 64'd1602731392, - 64'd942898944, - 64'd85956040, 64'd2398431739904, - 64'd1246460379136, 64'd136082161664, - 64'd585242, - 64'd988419008, - 64'd63059292, 64'd1787946991616, - 64'd1193769959424, 64'd146118590464, - 64'd1711474816, - 64'd1007434432, - 64'd39404984, 64'd1206294151168, - 64'd1131288723456, 64'd154783744000, - 64'd3505195520, - 64'd998888256, - 64'd15540209, 64'd658126929920, - 64'd1059999121408, 64'd161962950656, - 64'd5355531264, - 64'd962230336, 64'd7985572, 64'd147584860160, - 64'd980973191168, 64'd167563788288, - 64'd7235233792, - 64'd897425664, 64'd30631536, - 64'd321747517440, - 64'd895356567552, 64'd171517083648, - 64'd9116474368, - 64'd804953536, 64'd51876124, - 64'd746873421824, - 64'd804351574016, 64'd173777698816, - 64'd10971301888, - 64'd685797120, 64'd71227096, - 64'd1125407784960, - 64'd709200117760, 64'd174324940800, - 64'd12772102144, - 64'd541424320, 64'd88230856, - 64'd1455593095168, - 64'd611166257152, 64'd173162430464, - 64'd14492036096, - 64'd373759840, 64'd102480848, - 64'd1736305147904, - 64'd511518310400, 64'd170317807616, - 64'd16105472000, - 64'd185149968, 64'd113624944, - 64'd1967051767808, - 64'd411512045568, 64'd165841993728, - 64'd17588391936, 64'd21680196, 64'd121371688, - 64'd2147962060800, - 64'd312373608448, 64'd159808061440, - 64'd18918752256, 64'd243675424, 64'd125495320, - 64'd2279767277568, - 64'd215283679232, 64'd152309841920, - 64'd20076832768, 64'd477504352, 64'd125839424, - 64'd2363774205952, - 64'd121362456576, 64'd143460270080, - 64'd21045526528, 64'd719617600, 64'd122319368, - 64'd2401832534016, - 64'd31655704576, 64'd133389426688, - 64'd21810583552, 64'd966309248, 64'd114923288, - 64'd2396292644864, 64'd52877688832, 64'd122242334720, - 64'd22360815616, 64'd1213779968, 64'd103711792, - 64'd2349961052160, 64'd131376717824, 64'd110176616448, - 64'd22688249856, 64'd1458201344, 64'd88816312, - 64'd2266047971328, 64'd203087642624, 64'd97359986688, - 64'd22788214784, 64'd1695780224, 64'd70436248, - 64'd2148112007168, 64'd267371610112, 64'd83967647744, - 64'd22659383296, 64'd1922820864, 64'd48834932, - 64'd2000001302528, 64'd323710386176, 64'd70179553280, - 64'd22303770624, 64'd2135785856, 64'd24334446, - 64'd1825792065536, 64'd371710427136, 64'd56177754112, - 64'd21726658560, 64'd2331352832, - 64'd2690432, - 64'd1629725917184, 64'd411104739328, 64'd42143707136, - 64'd20936484864, 64'd2506467584, - 64'd31819196, - 64'd1416145666048, 64'd441753305088, 64'd28255617024, - 64'd19944681472, 64'd2658391808, - 64'd62593268, - 64'd1189433311232, 64'd463641182208, 64'd14685937664, - 64'd18765465600, 64'd2784744704, - 64'd94524208, - 64'd953947455488, 64'd476875259904, 64'd1598967424, - 64'd17415593984, 64'd2883539968, - 64'd127102344, - 64'd713963732992, 64'd481679081472, - 64'd10851364864, - 64'd15914071040, 64'd2953212672, - 64'd159805664, - 64'd473618382848, 64'd478386192384, - 64'd22523527168, - 64'd14281843712, 64'd2992642560, - 64'd192108752, - 64'd236854951936, 64'd467432079360, - 64'd33290172416, - 64'd12541457408, 64'd3001166848, - 64'd223491792, - 64'd7375633408, 64'd449344864256, - 64'd43039690752, - 64'd10716692480, 64'd2978587648, - 64'd253449152, 64'd211402358784, 64'd424734720000, - 64'd51677474816, - 64'd8832199680, 64'd2925170688, - 64'd281497824, 64'd416385105920, 64'd394282631168, - 64'd59126919168, - 64'd6913111040, 64'd2841636352, - 64'd307185344, 64'd604834299904, 64'd358728204288, - 64'd65330122752, - 64'd4984665088, 64'd2729145344, - 64'd330096832, 64'd774393626624, 64'd318857084928, - 64'd70248292352, - 64'd3071826176, 64'd2589274368, - 64'd349861728, 64'd923108311040, 64'd275487981568, - 64'd73861857280, - 64'd1198920320, 64'd2423989248, - 64'd366159488, 64'd1049438388224, 64'd229459607552, - 64'd76170289152, 64'd610715712, 64'd2235608832, - 64'd378724192, 64'd1152265617408, 64'd181617623040, - 64'd77191618560, 64'd2335062272, 64'd2026766848, - 64'd387348576, 64'd1230893875200, 64'd132802002944, - 64'd76961751040, 64'd3953719296, 64'd1800367104, - 64'd391886816, 64'd1285042470912, 64'd83834642432, - 64'd75533426688, 64'd5448179200, 64'd1559536128, - 64'd392256224, 64'd1314835398656, 64'd35507761152, - 64'd72975056896, 64'd6802064896, 64'd1307572608, - 64'd388438080, 64'd1320782528512, - 64'd11426966528, - 64'd69369282560, 64'd8001329664, 64'd1047895744, - 64'd380477152, 64'd1303757717504, - 64'd56268361728, - 64'd64811388928, 64'd9034421248, 64'd783991424, - 64'd368480608, 64'd1264970498048, - 64'd98374631424, - 64'd59407527936, 64'd9892401152, 64'd519358848, - 64'd352615392, 64'd1205935144960, - 64'd137171091456, - 64'd53272883200, 64'd10569023488, 64'd257457856, - 64'd333105184, 64'd1128434892800, - 64'd172156633088, - 64'd46529683456, 64'd11060770816, 64'd1657454, - 64'd310226112, 64'd1034484449280, - 64'd202908925952, - 64'd39305191424, 64'd11366848512, - 64'd244813248, - 64'd284301984, 64'd926288642048, - 64'd229088198656, - 64'd31729670144, 64'd11489137664, - 64'd478911104, - 64'd255698624, 64'd806201393152, - 64'd250439663616, - 64'd23934330880, 64'd11432105984, - 64'd697821312, - 64'd224817712, 64'd676682203136, - 64'd266794663936, - 64'd16049348608, 64'd11202685952, - 64'd898995520, - 64'd192090192, 64'd540253749248, - 64'd278070296576, - 64'd8201921536, 64'd10810113024, - 64'd1080185216, - 64'd157969200, 64'd399458729984, - 64'd284267872256, - 64'd514441984, 64'd10265736192, - 64'd1239470080, - 64'd122922824, 64'd256818872320, - 64'd285470064640, 64'd6897218048, 64'd9582800896, - 64'd1375280000, - 64'd87426824, 64'd114794971136, - 64'd281836912640, 64'd13925275648, 64'd8776203264, - 64'd1486412288, - 64'd51957212, - 64'd24250464256, - 64'd273600643072, 64'd20471439360, 64'd7862229504, - 64'd1572042496, - 64'd16983010, - 64'd158087888896, - 64'd261059772416, 64'd26448130048, 64'd6858277888, - 64'd1631729024, 64'd17040736, - 64'd284652142592, - 64'd244572110848, 64'd31779500032, 64'd5782572032, - 64'd1665412224, 64'd49679640, - 64'd402070208512, - 64'd224547143680, 64'd36402253824, 64'd4653866496, - 64'd1673407104, 64'd80526208, - 64'd508685058048, - 64'd201437888512, 64'd40266248192, 64'd3491151104, - 64'd1656391296, 64'd109205552, - 64'd603075248128, - 64'd175732293632, 64'd43334860800, 64'd2313361664, - 64'd1615386752, 64'd135380480, - 64'd684070141952, - 64'd147944243200, 64'd45585170432, 64'd1139094016, - 64'd1551737088, 64'd158755888, - 64'd750760820736, - 64'd118604644352, 64'd47007887360, - 64'd13666156, - 64'd1467081088, 64'd179082544, - 64'd802506014720, - 64'd88252309504, 64'd47607111680, - 64'd1127799296, - 64'd1363320832, 64'd196159872, - 64'd838934003712, - 64'd57425080320, 64'd47399833600, - 64'd2187287808, - 64'd1242587520, 64'd209838160, - 64'd859940061184, - 64'd26651252736, 64'd46415323136, - 64'd3177429760, - 64'd1107204736, 64'd220019792, - 64'd865679441920, 64'd3558628352, 64'd44694278144, - 64'd4085026560, - 64'd959648448, 64'd226659696, - 64'd856556503040, 64'd32719437824, 64'd42287857664, - 64'd4898542080, - 64'd802507008, 64'd229765008, - 64'd833210482688, 64'd60378497024, 64'd39256571904, - 64'd5608235008, - 64'd638439104, 64'd229393904, - 64'd796497477632, 64'd86121881600, 64'd35669041152, - 64'd6206257664, - 64'd470132416, 64'd225653632, - 64'd747469733888, 64'd109579927552, 64'd31600689152, - 64'd6686722048, - 64'd300262304, 64'd218697952, - 64'd687352250368, 64'd130431860736, 64'd27132338176, - 64'd7045738496, - 64'd131451952, 64'd208723776, - 64'd617517285376, 64'd148409516032, 64'd22348781568, - 64'd7281419776, 64'd33766012, 64'd195967312, - 64'd539457552384, 64'd163300114432, 64'd17337327616, - 64'd7393851392, 64'd192985360, 64'd180699632, - 64'd454757908480, 64'd174948057088, 64'd12186329088, - 64'd7385038848, 64'd343959488, 64'd163221824, - 64'd365066518528, 64'd183255728128, 64'd6983767040, - 64'd7258820096, 64'd484631296, 64'd143859824, - 64'd272065822720, 64'd188183445504, 64'd1815849472, - 64'd7020755456, 64'd613159616, 64'd122958880, - 64'd177443848192, 64'd189748363264, - 64'd3234301184, - 64'd6677993984, 64'd727941376, 64'd100877936, - 64'd82866216960, 64'd188022505472, - 64'd8087886336, - 64'd6239116800, 64'd827629760, 64'd77983912, 64'd10050632704, 64'd183130112000, - 64'd12671563776, - 64'd5713961984, 64'd911148096, 64'd54645936, 64'd99764699136, 64'd175244050432, - 64'd16918459392, - 64'd5113438208, 64'd977698944, 64'd31229768, 64'd184831721472, 64'd164581588992, - 64'd20769056768, - 64'd4449323008, 64'd1026768832, 64'd8092306, 64'd263926185984, 64'd151399677952, - 64'd24171935744, - 64'd3734053376, 64'd1058128640, - 64'd14423572, 64'd335859875840, 64'd135989600256, - 64'd27084365824, - 64'd2980513792, 64'd1071829056, - 64'd35993872, 64'd399597600768, 64'd118671261696, - 64'd29472751616, - 64'd2201821440, 64'd1068192768, - 64'd56317924, 64'd454270091264, 64'd99787186176, - 64'd31312910336, - 64'd1411112448, 64'd1047801408, - 64'd75122352, 64'd499183616000, 64'd79696314368, - 64'd32590198784, - 64'd621336384, 64'd1011480128, - 64'd92164568, 64'd533826732032, 64'd58767691776, - 64'd33299482624, 64'd154943552, 64'd960277760, - 64'd107235656, 64'd557873823744, 64'd37374169088, - 64'd33444954112, 64'd905737024, 64'd895444608, - 64'd120162680, 64'd571185233920, 64'd15886231552, - 64'd33039812608, 64'd1619800192, 64'd818407360, - 64'd130810440, 64'd573804773376, - 64'd5333987328, - 64'd32105801728, 64'd2286791936, 64'd730742464, - 64'd139082496, 64'd565953953792, - 64'd25938384896, - 64'd30672625664, 64'd2897413120, 64'd634146880, - 64'd144921664, 64'd548023926784, - 64'd45598187520, - 64'd28777254912, 64'd3443524096, 64'd530409024, - 64'd148309872, 64'd520564146176, - 64'd64008802304, - 64'd26463137792, 64'd3918241280, 64'd421377696, - 64'd149267344, 64'd484269522944, - 64'd80894140416, - 64'd23779321856, 64'd4316012544, 64'd308932032, - 64'd147851344, 64'd439965057024, - 64'd96010354688, - 64'd20779517952, 64'd4632668160, 64'd194951008, - 64'd144154208, 64'd388588961792, - 64'd109148995584, - 64'd17521113088, 64'd4865448448, 64'd81284144, - 64'd138301056, 64'd331174313984, - 64'd120139448320, - 64'd14064135168, 64'd5013009408, - 64'd30276684, - 64'd130446984, 64'd268829605888, - 64'd128850771968, - 64'd10470236160, 64'd5075404800, - 64'd138023792, - 64'd120773768, 64'd202718658560, - 64'd135192780800, - 64'd6801641472, 64'd5054048768, - 64'd240358176, - 64'd109486384, 64'd134040117248, - 64'd139116445696, - 64'd3120139008, 64'd4951653888, - 64'd335811680, - 64'd96809216, 64'd64006848512, - 64'd140613697536, 64'd513904608, 64'd4772154368, - 64'd423066464, - 64'd82981984, - 64'd6174270464, - 64'd139716444160, 64'd4042478336, 64'd4520609792, - 64'd500971680, - 64'd68255632, - 64'd75322032128, - 64'd136495087616, 64'd7410798592, 64'd4203092992, - 64'd568556992, - 64'd52888100, - 64'd142299611136, - 64'd131056402432, 64'd10568109056, 64'd3826567936, - 64'd625043008, - 64'd37140108, - 64'd206032109568, - 64'd123540840448, 64'd13468387328, 64'd3398753024, - 64'd669848256, - 64'd21271010, - 64'd265522659328, - 64'd114119467008, 64'd16070970368, 64'd2927977984, - 64'd702593088, - 64'd5534769, - 64'd319866830848, - 64'd102990364672, 64'd18341064704, 64'd2423034880, - 64'd723099968, 64'd9823876, - 64'd368265166848, - 64'd90374766592, 64'd20250150912, 64'd1893024640, - 64'd731391104, 64'd24572992, - 64'd410033782784, - 64'd76512894976, 64'd21776293888, 64'd1347204352, - 64'd727682368, 64'd38496744, - 64'd444612771840, - 64'd61659594752, 64'd22904309760, 64'd794834368, - 64'd712374656, 64'd51398352, - 64'd471572283392, - 64'd46079827968, 64'd23625850880, 64'd245030640, - 64'd686042560, 64'd63102660, - 64'd490616586240, - 64'd30044149760, 64'd23939354624, - 64'd293377280, - 64'd649420608, 64'd73458312, - 64'd501585739776, - 64'd13824169984, 64'd23849902080, - 64'd811979904, - 64'd603387136, 64'd82339488, - 64'd504454807552, 64'd2311850496, 64'd23368964096, - 64'd1302911104, - 64'd548946496, 64'd89647192, - 64'd499331366912, 64'd18103277568, 64'd22514049024, - 64'd1758959872, - 64'd487209728, 64'd95310104, - 64'd486450528256, 64'd33301121024, 64'd21308276736, - 64'd2173667840, - 64'd419373920, 64'd99284920, - 64'd466168217600, 64'd47671787520, 64'd19779858432, - 64'd2541413888, - 64'd346700928, 64'd101556320, - 64'd438952525824, 64'd61000474624, 64'd17961517056, - 64'd2857481216, - 64'd270495520, 64'd102136416, - 64'd405373714432, 64'd73094193152, 64'd15889840128, - 64'd3118109184, - 64'd192083456, 64'd101063864, - 64'd366092419072, 64'd83784359936, 64'd13604604928, - 64'd3320529664, - 64'd112789768, 64'd98402488, - 64'd321847099392, 64'd92928925696, 64'd11148049408, - 64'd3462983936, - 64'd33917672, 64'd94239632, - 64'd273440227328, 64'd100414029824, 64'd8564135936, - 64'd3544725760, 64'd43271628, 64'd88684120, - 64'd221723901952, 64'd106155171840, 64'd5897799168, - 64'd3566006272, 64'd117577960, 64'd81863952, - 64'd167584972800, 64'd110097866752, 64'd3194200576, - 64'd3528044544, 64'd187879696, 64'd73923784, - 64'd111929999360, 64'd112217784320, 64'd497996768, - 64'd3432982528, 64'd253149584, 64'd65022140, - 64'd55670218752, 64'd112520486912, - 64'd2147366144, - 64'd3283827200, 64'd312468704, 64'd55328580, 64'd293226432, 64'd111040561152, - 64'd4700319744, - 64'd3084379648, 64'd365038144, 64'd45020656, 64'd55083495424, 64'd107840413696, - 64'd7121794560, - 64'd2839154688, 64'd410188800, 64'd34280916, 64'd107861565440, 64'd103008600064, - 64'd9375787008, - 64'd2553288192, 64'd447388512, 64'd23293848, 64'd157838802944, 64'd96657784832, - 64'd11429858304, - 64'd2232440832, 64'd476246976, 64'd12242892, 64'd204288475136, 64'd88922374144, - 64'd13255571456, - 64'd1882692224, 64'd496518336, 64'd1307557, 64'd246555901952, 64'd79955836928, - 64'd14828847104, - 64'd1510434048, 64'd508101280, - 64'd9339338, 64'd284067299328, 64'd69927788544, - 64'd16130240512, - 64'd1122258432, 64'd511036928, - 64'd19534240, 64'd316337160192, 64'd59020926976, - 64'd17145144320, - 64'd724847744, 64'd505504416, - 64'd29125226, 64'd342973808640, 64'd47427776512, - 64'd17863899136, - 64'd324865088, 64'd491814400, - 64'd37974108, 64'd363683708928, 64'd35347369984, - 64'd18281832448, 64'd71152392, 64'd470400736, - 64'd45958284, 64'd378273693696, 64'd22981933056, - 64'd18399207424, 64'd456894976, 64'd441810336, - 64'd52972284, 64'd386651848704, 64'd10533573632, - 64'd18221096960, 64'd826375808, 64'd406691392, - 64'd58928988, 64'd388826595328, - 64'd1798948096, - 64'd17757192192, 64'd1174018944, 64'd365780480, - 64'd63760556, 64'd384904298496, - 64'd13823309824, - 64'd17021529088, 64'd1494738304, 64'd319888416, - 64'd67418992, 64'd375085203456, - 64'd25356541952, - 64'd16032155648, 64'd1784006784, 64'd269885376, - 64'd69876376, 64'd359658192896, - 64'd36227723264, - 64'd14810752000, 64'd2037915392, 64'd216685360, - 64'd71124832, 64'd338994003968, - 64'd46280421376, - 64'd13382192128, 64'd2253219584, 64'd161230592, - 64'd71176072, 64'd313537560576, - 64'd55374839808, - 64'd11774067712, 64'd2427375104, 64'd104475496, - 64'd70060744, 64'd283799191552, - 64'd63389650944, - 64'd10016183296, 64'd2558562304, 64'd47371200, - 64'd67827424, 64'd250344865792, - 64'd70223495168, - 64'd8140022272, 64'd2645694720, - 64'd9149640, - 64'd64541392, 64'd213786034176, - 64'd75796103168, - 64'd6178208256, 64'd2688421120, - 64'd64187332, - 64'd60283132, 64'd174768832512, - 64'd80049086464, - 64'd4163952384, 64'd2687111168, - 64'd116888728, - 64'd55146664, 64'd133963022336, - 64'd82946351104, - 64'd2130511360, 64'd2642831616, - 64'd166459696, - 64'd49237692, 64'd92050849792, - 64'd84474118144, - 64'd110653576, 64'd2557312768, - 64'd212176416, - 64'd42671612, 64'd49715904512, - 64'd84640620544, 64'd1863850752, 64'd2432903936, - 64'd253395088, - 64'd35571408, 64'd7632287232, - 64'd83475464192, 64'd3762712832, 64'd2272520192, - 64'd289560384, - 64'd28065490, - 64'd33545834496, - 64'd81028612096, 64'd5557572608, 64'd2079582848, - 64'd320211968, - 64'd20285500, - 64'd73194119168, - 64'd77369139200, 64'd7222403072, 64'd1857950848, - 64'd344989568, - 64'd12364129, - 64'd110727217152, - 64'd72583659520, 64'd8733871104, 64'd1611849088, - 64'd363636256, - 64'd4432954, - 64'd145607098368, - 64'd66774532096, 64'd10071640064, 64'd1345791744, - 64'd375999936, 64'd3379635, - 64'd177350426624, - 64'd60057858048, 64'd11218626560, 64'd1064502912, - 64'd382033088, 64'd10950404, - 64'd205534920704, - 64'd52561313792, 64'd12161187840, 64'd772835904, - 64'd381791072, 64'd18163128, - 64'd229804539904, - 64'd44421840896, 64'd12889261056, 64'd475692544, - 64'd375428544, 64'd24910266, - 64'd249873547264, - 64'd35783254016, 64'd13396432896, 64'd177943536, - 64'd363194560, 64'd31094466, - 64'd265529311232, - 64'd26793799680, 64'd13679954944, - 64'd115648360, - 64'd345426240, 64'd36629864, - 64'd276633911296, - 64'd17603684352, 64'd13740696576, - 64'd400501952, - 64'd322541184, 64'd41443168, - 64'd283124531200, - 64'd8362662400, 64'd13583045632, - 64'd672286208, - 64'd295028768, 64'd45474524, - 64'd285012590592, 64'd782341184, 64'd13214753792, - 64'd926983424, - 64'd263440544, 64'd48678116, - 64'd282381877248, 64'd9689481216, 64'd12646726656, - 64'd1160945536, - 64'd228379888, 64'd51022572, - 64'd275385253888, 64'd18224119808, 64'd11892779008, - 64'd1370943232, - 64'd190491040, 64'd52491072, - 64'd264240807936, 64'd26260789248, 64'd10969340928, - 64'd1554207488, - 64'd150447840, 64'd53081284, - 64'd249226625024, 64'd33684951040, 64'd9895136256, - 64'd1708462336, - 64'd108942160, 64'd52805020, - 64'd230675021824, 64'd40394547200, 64'd8690825216, - 64'd1831949184, - 64'd66672452, 64'd51687692, - 64'd208965959680, 64'd46301310976, 64'd7378630656, - 64'd1923442048, - 64'd24332392, 64'd49767576, - 64'd184519835648, 64'd51331833856, 64'd5981947904, - 64'd1982254208, 64'd17400088, 64'd47094876, - 64'd157789880320, 64'd55428366336, 64'd4524942848, - 64'd2008235904, 64'd57873236, 64'd43730612, - 64'd129254154240, 64'd58549334016, 64'd3032150016, - 64'd2001763840, 64'd96471240, 64'd39745388, - 64'd99407421440, 64'd60669616128, 64'd1528072832, - 64'd1963721984, 64'd132623208, 64'd35218024, - 64'd68752859136, 64'd61780545536, 64'd36796504, - 64'd1895475328, 64'd165811136, 64'd30234082, - 64'd37793939456, 64'd61889617920, - 64'd1418385152, - 64'd1798836224, 64'd195576944, 64'd24884336, - 64'd7026437632, 64'd61020004352, - 64'd2815320320, - 64'd1676024704, 64'd221528240, 64'd19263196, 64'd23069216768, 64'd59209773056, - 64'd4133322240, - 64'd1529623168, 64'd243343024, 64'd13467098, 64'd52035162112, 64'd56510943232, - 64'd5353462784, - 64'd1362526464, 64'd260773104, 64'd7592925, 64'd79442788352, 64'd52988293120, - 64'd6458829824, - 64'd1177887744, 64'd273646208, 64'd1736438, 64'd104898797568, 64'd48718045184, - 64'd7434744832, - 64'd979062912, 64'd281866912, - 64'd4009222, 64'd128050544640, 64'd43786350592, - 64'd8268942848, - 64'd769551040, 64'd285416224, - 64'd9554955, 64'd148590624768, 64'd38287704064, - 64'd8951707648, - 64'd552936192, 64'd284350048, - 64'd14817033, 64'd166260588544, 64'd32323217408, - 64'd9475960832, - 64'd332827776, 64'd278796512, - 64'd19718296, 64'd180853850112, 64'd25998870528, - 64'd9837315072, - 64'd112802824, 64'd268952064, - 64'd24189226, 64'd192217645056, 64'd19423698944, - 64'd10034070528, 64'd103650368, 64'd255076688, - 64'd28168872, 64'd200254128128, 64'd12708000768, - 64'd10067181568, 64'd313185376, 64'd237488272, - 64'd31605606, 64'd204920520704, 64'd5961550848, - 64'd9940171776, 64'd512647424, 64'd216556032, - 64'd34457716, 64'd206228488192, - 64'd708124480, - 64'd9659018240, 64'd699118848, 64'd192693456, - 64'd36693844, 64'd204242501632, - 64'd7197395456, - 64'd9231992832, 64'd869959680, 64'd166350592, - 64'd38293204, 64'd199077560320, - 64'd13408075776, - 64'd8669478912, 64'd1022842816, 64'd138005968, - 64'd39245684, 64'd190896128000, - 64'd19248842752, - 64'd7983748096, 64'd1155783296, 64'd108158320, - 64'd39551716, 64'd179904282624, - 64'd24636518400, - 64'd7188726272, 64'd1267161216, 64'd77318152, - 64'd39222040, 64'd166347489280, - 64'd29497176064, - 64'd6299724288, 64'd1355739264, 64'd45999272, - 64'd38277248, 64'd150505635840, - 64'd33767094272, - 64'd5333166592, 64'd1420672000, 64'd14710599, - 64'd36747244, 64'd132687716352, - 64'd37393506304, - 64'd4306299904, 64'd1461510272, - 64'd16051860, - 64'd34670516, 64'd113226309632, - 64'd40335167488, - 64'd3236899328, 64'd1478198528, - 64'd45812568, - 64'd32093330, 64'd92471631872, - 64'd42562719744, - 64'd2142974848, 64'd1471065856, - 64'd74123520, - 64'd29068780, 64'd70785564672, - 64'd44058857472, - 64'd1042477568, 64'd1440811392, - 64'd100570712, - 64'd25655798, 64'd48535621632, - 64'd44818313216, 64'd46982476, 64'd1388484224, - 64'd124779864, - 64'd21918058, 64'd26089003008, - 64'd44847632384, 64'd1108407680, 64'd1315457664, - 64'd146421424, - 64'd17922850, 64'd3806748672, - 64'd44164767744, 64'd2125667584, 64'd1223400064, - 64'd165214688, - 64'd13739916, - 64'd17961811968, - 64'd42798526464, 64'd3083733504, 64'd1114240512, - 64'd180931088, - 64'd9440287, - 64'd38884319232, - 64'd40787836928, 64'd3968889600, 64'd990132288, - 64'd193396528, - 64'd5095112, - 64'd58650222592, - 64'd38180864000, 64'd4768918016, 64'd853412352, - 64'd202492816, - 64'd774528, - 64'd76975161344, - 64'd35034038272, 64'd5473255936, 64'd706560576, - 64'd208158176, 64'd3453433, - 64'd93604839424, - 64'd31410925568, 64'd6073121280, 64'd552156160, - 64'd210386848, 64'd7523876, - 64'd108318269440, - 64'd27381069824, 64'd6561609728, 64'd392834496, - 64'd209227760, 64'd11375996, - 64'd120930476032, - 64'd23018717184, 64'd6933754880, 64'd231244032, - 64'd204782480, 64'd14953949, - 64'd131294502912, - 64'd18401529856, 64'd7186563072, 64'd70003600, - 64'd197202240, 64'd18207614, - 64'd139302813696, - 64'd13609263104, 64'd7319006720, - 64'd88338248, - 64'd186684336, 64'd21093252, - 64'd144888004608, - 64'd8722452480, 64'd7331995648, - 64'd241342064, - 64'd173467872, 64'd23574048, - 64'd148022853632, - 64'd3821109760, 64'd7228313600, - 64'd386713472, - 64'd157828880, 64'd25620520, - 64'd148719747072, 64'd1016530176, 64'd7012526592, - 64'd522336128, - 64'd140075104, 64'd27210812, - 64'd147029508096, 64'd5715210240, 64'd6690865664, - 64'd646300800, - 64'd120540240, 64'd28330850, - 64'd143039594496, 64'd10203770880, 64'd6271088640, - 64'd756930624, - 64'd99578080, 64'd28974380, - 64'd136871796736, 64'd14416177152, 64'd5762317312, - 64'd852802112, - 64'd77556320, 64'd29142874, - 64'd128679477248, 64'd18292439040, 64'd5174857728, - 64'd932761088, - 64'd54850424, 64'd28845310, - 64'd118644285440, 64'd21779417088, 64'd4520009728, - 64'd995934912, - 64'd31837438, 64'd28097850, - 64'd106972594176, 64'd24831485952, 64'd3809860352, - 64'd1041738880, - 64'd8889991, 64'd26923408, - 64'd93891592192, 64'd27411083264, 64'd3057072896, - 64'd1069878528, 64'd13629545, 64'd25351112, - 64'd79645155328, 64'd29489094656, 64'd2274671616, - 64'd1080347136, 64'd35374540, 64'd23415698, - 64'd64489545728, 64'd31045109760, 64'd1475826304, - 64'd1073418880, 64'd56019228, 64'd21156812, - 64'd48689025024, 64'd32067528704, 64'd673638400, - 64'd1049637120, 64'd75263368, 64'd18618256, - 64'd32511469568, 64'd32553523200, - 64'd119064600, - 64'd1009799232, 64'd92836392, 64'd15847203, - 64'd16223992832, 64'd32508864512, - 64'd889926592, - 64'd954937920, 64'd108500936, 64'd12893350, - 64'd88746856, 64'd31947616256, - 64'd1627247104, - 64'd886298624, 64'd122055824, 64'd9808074, 64'd15641138176, 64'd30891702272, - 64'd2320150784, - 64'd805314432, 64'd133338360, 64'd6643568, 64'd30725345280, 64'd29370359808, - 64'd2958740480, - 64'd713579008, 64'd142225952, 64'd3452002, 64'd44939878400, 64'd27419498496, - 64'd3534228480, - 64'd612817024, 64'd148637040, 64'd284680, 64'd58080198656, 64'd25080952832, - 64'd4039049984, - 64'd504853440, 64'd152531456, - 64'd2808740, 64'd69964013568, 64'd22401675264, - 64'd4466952192, - 64'd391582240, 64'd153909936, - 64'd5781004, 64'd80433602560, 64'd19432865792, - 64'd4813060608, - 64'd274934528, 64'd152813168, - 64'd8587947, 64'd89357697024, 64'd16229040128, - 64'd5073922560, - 64'd156846864, 64'd149320128, - 64'd11189123, 64'd96632946688, 64'd12847086592, - 64'd5247527424, - 64'd39230476, 64'd143545872, - 64'd13548353, 64'd102184812544, 64'd9345304576, - 64'd5333300736, 64'd76058528, 64'd135638800, - 64'd15634194, 64'd105968074752, 64'd5782438912, - 64'd5332078080, 64'd187247280, 64'd125777552, - 64'd17420324, 64'd107966783488, 64'd2216733952, - 64'd5246058496, 64'd292672224, 64'd114167280, - 64'd18885832, 64'd108193816576, - 64'd1294978432, - 64'd5078732800, 64'd390802848, 64'd101035864, - 64'd20015412, 64'd106689912832, - 64'd4698147328, - 64'd4834797056, 64'd480262688, 64'd86629656, - 64'd20799476, 64'd103522353152, - 64'd7941314048, - 64'd4520049152, 64'd559847360, 64'd71209128, - 64'd21234158, 64'd98783232000, - 64'd10976852992, - 64'd4141266432, 64'd628539328, 64'd55044372, - 64'd21321234, 64'd92587327488, - 64'd13761633280, - 64'd3706075648, 64'd685519616, 64'd38410596, - 64'd21067960, 64'd85069766656, - 64'd16257591296, - 64'd3222810112, 64'd730175616, 64'd21583592, - 64'd20486812, 64'd76383322112, - 64'd18432212992, - 64'd2700358656, 64'd762106048, 64'd4835369, - 64'd19595166, 64'd66695573504, - 64'd20258908160, - 64'd2148011520, 64'd781121600, - 64'd11570094, - 64'd18414896, 64'd56185835520, - 64'd21717288960, - 64'd1575302784, 64'd787243072, - 64'd27380832, - 64'd16971916, 64'd45042040832, - 64'd22793334784, - 64'd991851136, 64'd780695552, - 64'd42360600, - 64'd15295670, 64'd33457522688, - 64'd23479463936, - 64'd407206720, 64'd761899904, - 64'd56292244, - 64'd13418574, 64'd21627799552, - 64'd23774482432, 64'd169300192, 64'd731461184, - 64'd68980656, - 64'd11375428, 64'd9747416064, - 64'd23683454976, 64'd728701632, 64'd690154240, - 64'd80255344, - 64'd9202805, - 64'd1993129344, - 64'd23217463296, 64'd1262525568, 64'd638907456, - 64'd89972536, - 64'd6938424, - 64'd13410318336, - 64'd22393276416, 64'd1762918144, 64'd578783936, - 64'd98016768, - 64'd4620524, - 64'd24330354688, - 64'd21232945152, 64'd2222753536, 64'd510961472, - 64'd104302040, - 64'd2287246, - 64'd34591690752, - 64'd19763324928, 64'd2635728128, 64'd436710720, - 64'd108772432, 64'd23980, - 64'd44047294464, - 64'd18015514624, 64'd2996441856, 64'd357372896, - 64'd111402280, 64'd2276999, - 64'd52566618112, - 64'd16024272896, 64'd3300460032, 64'd274336512, - 64'd112195776, 64'd4437484, - 64'd60037275648, - 64'd13827361792, 64'd3544360448, 64'd189014320, - 64'd111186200, 64'd6473431, - 64'd66366373888, - 64'd11464875008, 64'd3725762560, 64'd102820136, - 64'd108434648, 64'd8355611, - 64'd71481499648, - 64'd8978542592, 64'd3843339264, 64'd17146324, - 64'd104028384, 64'd10057966, - 64'd75331379200, - 64'd6411025408, 64'd3896812032, - 64'd66657732, - 64'd98078776, 64'd11557943, - 64'd77886144512, - 64'd3805214208, 64'd3886928128, - 64'd147306064, - 64'd90718944, 64'd12836766, - 64'd79137292288, - 64'd1203540608, 64'd3815425280, - 64'd223594944, - 64'd82101112, 64'd13879640, - 64'd79097274368, 64'd1352686720, 64'd3684976896, - 64'd294420000, - 64'd72393696, 64'd14675887, - 64'd77798785024, 64'd3823910656, 64'd3499128064, - 64'd358791296, - 64'd61778220, 64'd15219014, - 64'd75293745152, 64'd6172911616, 64'd3262216448, - 64'd415846208, - 64'd50446116, 64'd15506713, - 64'd71651991552, 64'd8365341184, 64'd2979283968, - 64'd464859936, - 64'd38595436, 64'd15540788, - 64'd66959687680, 64'd10370196480, 64'd2655979008, - 64'd505253664, - 64'd26427528, 64'd15327032, - 64'd61317615616, 64'd12160233472, 64'd2298451200, - 64'd536600032, - 64'd14143770, 64'd14875031, - 64'd54839140352, 64'd13712301056, 64'd1913241984, - 64'd558626304, - 64'd1942347, 64'd14197915, - 64'd47648133120, 64'd15007612928, 64'd1507169536, - 64'd571214592, 64'd9984802, 64'd13312069, - 64'd39876722688, 64'd16031933440, 64'd1087214208, - 64'd574400256, 64'd21454888, 64'd12236782, - 64'd31662987264, 64'd16775695360, 64'd660403712, - 64'd568367104, 64'd32296946, 64'd10993875, - 64'd23148623872, 64'd17234030592, 64'd233699392, - 64'd553441088, 64'd42354264, 64'd9607290, - 64'd14476587008, 64'd17406736384, - 64'd186112288, - 64'd530081408, 64'd51486508, 64'd8102654, - 64'd5788791296, 64'd17298159616, - 64'd592523456, - 64'd498869920, 64'd59571556, 64'd6506830, 64'd2776121088, 64'd16917010432, - 64'd979401536, - 64'd460498944, 64'd66506984, 64'd4847465, 64'd11084907520, 64'd16276123648, - 64'd1341077248, - 64'd415757280, 64'd72211192, 64'd3152522, 64'd19011708928, 64'd15392145408, - 64'd1672423168, - 64'd365515520, 64'd76624208, 64'd1449835, 64'd26439870464, 64'd14285174784, - 64'd1968922496, - 64'd310709952, 64'd79708064, - 64'd233334, 64'd33263562752, 64'd12978362368, - 64'd2226724608, - 64'd252326112, 64'd81446888, - 64'd1870714, 64'd39389204480, 64'd11497459712, - 64'd2442690560, - 64'd191381936, 64'd81846584, - 64'd3437414, 64'd44736643072, 64'd9870348288, - 64'd2614424576, - 64'd128910704, 64'd80934216, - 64'd4910289};
	localparam logic signed[63:0] hb[0:1799] = {64'd11671469817856, 64'd68906754048, - 64'd75389681664, - 64'd632993600, 64'd1232912256, 64'd13692950, 64'd11602687426560, 64'd205972455424, - 64'd73580404736, - 64'd1884879744, 64'd1207679872, 64'd40773932, 64'd11465870278656, 64'd340804698112, - 64'd69988712448, - 64'd3094723328, 64'd1157783296, 64'd66948644, 64'd11262497914880, 64'd471947444224, - 64'd64667860992, - 64'd4235354880, 64'd1084343936, 64'd91640440, 64'd10994772344832, 64'd597993521152, - 64'd57696690176, - 64'd5280870912, 64'd989008640, 64'd114312056, 64'd10665578201088, 64'd717603078144, - 64'd49178345472, - 64'd6207100416, 64'd873910592, 64'd134478512, 64'd10278451281920, 64'd829521199104, - 64'd39238668288, - 64'd6992039424, 64'd741620736, 64'd151718128, 64'd9837531365376, 64'd932594057216, - 64'd28024207360, - 64'd7616239104, 64'd595090240, 64'd165681392, 64'd9347505586176, 64'd1025783496704, - 64'd15699915776, - 64'd8063150592, 64'd437586208, 64'd176098000, 64'd8813547618304, 64'd1108180467712, - 64'd2446590720, - 64'd8319411200, 64'd272621824, 64'd182781520, 64'd8241252663296, 64'd1179015708672, 64'd11541940224, - 64'd8375070720, 64'd103882200, 64'd185632240, 64'd7636563001344, 64'd1237668986880, 64'd26061805568, - 64'd8223759872, - 64'd64851640, 64'd184637792, 64'd7005691969536, 64'd1283676045312, 64'd40902221824, - 64'd7862790656, - 64'd229779984, 64'd179871936, 64'd6355046367232, 64'd1316733190144, 64'd55848693760, - 64'd7293190144, - 64'd387160704, 64'd171491536, 64'd5691141521408, 64'd1336699518976, 64'd70686261248, - 64'd6519671296, - 64'd533383328, 64'd159731776, 64'd5020525789184, 64'd1343597314048, 64'd85202714624, - 64'd5550539264, - 64'd665039680, 64'd144899840, 64'd4349692739584, 64'd1337609420800, 64'd99191758848, - 64'd4397536256, - 64'd778989504, 64'd127367376, 64'd3685008015360, 64'd1319074791424, 64'd112455999488, - 64'd3075626240, - 64'd872420032, 64'd107561680, 64'd3032628592640, 64'd1288481931264, 64'd124809854976, - 64'd1602731392, - 64'd942898944, 64'd85956040, 64'd2398431739904, 64'd1246460379136, 64'd136082161664, 64'd585242, - 64'd988419008, 64'd63059292, 64'd1787946991616, 64'd1193769959424, 64'd146118590464, 64'd1711474816, - 64'd1007434432, 64'd39404984, 64'd1206294151168, 64'd1131288723456, 64'd154783744000, 64'd3505195520, - 64'd998888256, 64'd15540209, 64'd658126929920, 64'd1059999121408, 64'd161962950656, 64'd5355531264, - 64'd962230336, - 64'd7985572, 64'd147584860160, 64'd980973191168, 64'd167563788288, 64'd7235233792, - 64'd897425664, - 64'd30631536, - 64'd321747517440, 64'd895356567552, 64'd171517083648, 64'd9116474368, - 64'd804953536, - 64'd51876124, - 64'd746873421824, 64'd804351574016, 64'd173777698816, 64'd10971301888, - 64'd685797120, - 64'd71227096, - 64'd1125407784960, 64'd709200117760, 64'd174324940800, 64'd12772102144, - 64'd541424320, - 64'd88230856, - 64'd1455593095168, 64'd611166257152, 64'd173162430464, 64'd14492036096, - 64'd373759840, - 64'd102480848, - 64'd1736305147904, 64'd511518310400, 64'd170317807616, 64'd16105472000, - 64'd185149968, - 64'd113624944, - 64'd1967051767808, 64'd411512045568, 64'd165841993728, 64'd17588391936, 64'd21680196, - 64'd121371688, - 64'd2147962060800, 64'd312373608448, 64'd159808061440, 64'd18918752256, 64'd243675424, - 64'd125495320, - 64'd2279767277568, 64'd215283679232, 64'd152309841920, 64'd20076832768, 64'd477504352, - 64'd125839424, - 64'd2363774205952, 64'd121362456576, 64'd143460270080, 64'd21045526528, 64'd719617600, - 64'd122319368, - 64'd2401832534016, 64'd31655704576, 64'd133389426688, 64'd21810583552, 64'd966309248, - 64'd114923288, - 64'd2396292644864, - 64'd52877688832, 64'd122242334720, 64'd22360815616, 64'd1213779968, - 64'd103711792, - 64'd2349961052160, - 64'd131376717824, 64'd110176616448, 64'd22688249856, 64'd1458201344, - 64'd88816312, - 64'd2266047971328, - 64'd203087642624, 64'd97359986688, 64'd22788214784, 64'd1695780224, - 64'd70436248, - 64'd2148112007168, - 64'd267371610112, 64'd83967647744, 64'd22659383296, 64'd1922820864, - 64'd48834932, - 64'd2000001302528, - 64'd323710386176, 64'd70179553280, 64'd22303770624, 64'd2135785856, - 64'd24334446, - 64'd1825792065536, - 64'd371710427136, 64'd56177754112, 64'd21726658560, 64'd2331352832, 64'd2690432, - 64'd1629725917184, - 64'd411104739328, 64'd42143707136, 64'd20936484864, 64'd2506467584, 64'd31819196, - 64'd1416145666048, - 64'd441753305088, 64'd28255617024, 64'd19944681472, 64'd2658391808, 64'd62593268, - 64'd1189433311232, - 64'd463641182208, 64'd14685937664, 64'd18765465600, 64'd2784744704, 64'd94524208, - 64'd953947455488, - 64'd476875259904, 64'd1598967424, 64'd17415593984, 64'd2883539968, 64'd127102344, - 64'd713963732992, - 64'd481679081472, - 64'd10851364864, 64'd15914071040, 64'd2953212672, 64'd159805664, - 64'd473618382848, - 64'd478386192384, - 64'd22523527168, 64'd14281843712, 64'd2992642560, 64'd192108752, - 64'd236854951936, - 64'd467432079360, - 64'd33290172416, 64'd12541457408, 64'd3001166848, 64'd223491792, - 64'd7375633408, - 64'd449344864256, - 64'd43039690752, 64'd10716692480, 64'd2978587648, 64'd253449152, 64'd211402358784, - 64'd424734720000, - 64'd51677474816, 64'd8832199680, 64'd2925170688, 64'd281497824, 64'd416385105920, - 64'd394282631168, - 64'd59126919168, 64'd6913111040, 64'd2841636352, 64'd307185344, 64'd604834299904, - 64'd358728204288, - 64'd65330122752, 64'd4984665088, 64'd2729145344, 64'd330096832, 64'd774393626624, - 64'd318857084928, - 64'd70248292352, 64'd3071826176, 64'd2589274368, 64'd349861728, 64'd923108311040, - 64'd275487981568, - 64'd73861857280, 64'd1198920320, 64'd2423989248, 64'd366159488, 64'd1049438388224, - 64'd229459607552, - 64'd76170289152, - 64'd610715712, 64'd2235608832, 64'd378724192, 64'd1152265617408, - 64'd181617623040, - 64'd77191618560, - 64'd2335062272, 64'd2026766848, 64'd387348576, 64'd1230893875200, - 64'd132802002944, - 64'd76961751040, - 64'd3953719296, 64'd1800367104, 64'd391886816, 64'd1285042470912, - 64'd83834642432, - 64'd75533426688, - 64'd5448179200, 64'd1559536128, 64'd392256224, 64'd1314835398656, - 64'd35507761152, - 64'd72975056896, - 64'd6802064896, 64'd1307572608, 64'd388438080, 64'd1320782528512, 64'd11426966528, - 64'd69369282560, - 64'd8001329664, 64'd1047895744, 64'd380477152, 64'd1303757717504, 64'd56268361728, - 64'd64811388928, - 64'd9034421248, 64'd783991424, 64'd368480608, 64'd1264970498048, 64'd98374631424, - 64'd59407527936, - 64'd9892401152, 64'd519358848, 64'd352615392, 64'd1205935144960, 64'd137171091456, - 64'd53272883200, - 64'd10569023488, 64'd257457856, 64'd333105184, 64'd1128434892800, 64'd172156633088, - 64'd46529683456, - 64'd11060770816, 64'd1657454, 64'd310226112, 64'd1034484449280, 64'd202908925952, - 64'd39305191424, - 64'd11366848512, - 64'd244813248, 64'd284301984, 64'd926288642048, 64'd229088198656, - 64'd31729670144, - 64'd11489137664, - 64'd478911104, 64'd255698624, 64'd806201393152, 64'd250439663616, - 64'd23934330880, - 64'd11432105984, - 64'd697821312, 64'd224817712, 64'd676682203136, 64'd266794663936, - 64'd16049348608, - 64'd11202685952, - 64'd898995520, 64'd192090192, 64'd540253749248, 64'd278070296576, - 64'd8201921536, - 64'd10810113024, - 64'd1080185216, 64'd157969200, 64'd399458729984, 64'd284267872256, - 64'd514441984, - 64'd10265736192, - 64'd1239470080, 64'd122922824, 64'd256818872320, 64'd285470064640, 64'd6897218048, - 64'd9582800896, - 64'd1375280000, 64'd87426824, 64'd114794971136, 64'd281836912640, 64'd13925275648, - 64'd8776203264, - 64'd1486412288, 64'd51957212, - 64'd24250464256, 64'd273600643072, 64'd20471439360, - 64'd7862229504, - 64'd1572042496, 64'd16983010, - 64'd158087888896, 64'd261059772416, 64'd26448130048, - 64'd6858277888, - 64'd1631729024, - 64'd17040736, - 64'd284652142592, 64'd244572110848, 64'd31779500032, - 64'd5782572032, - 64'd1665412224, - 64'd49679640, - 64'd402070208512, 64'd224547143680, 64'd36402253824, - 64'd4653866496, - 64'd1673407104, - 64'd80526208, - 64'd508685058048, 64'd201437888512, 64'd40266248192, - 64'd3491151104, - 64'd1656391296, - 64'd109205552, - 64'd603075248128, 64'd175732293632, 64'd43334860800, - 64'd2313361664, - 64'd1615386752, - 64'd135380480, - 64'd684070141952, 64'd147944243200, 64'd45585170432, - 64'd1139094016, - 64'd1551737088, - 64'd158755888, - 64'd750760820736, 64'd118604644352, 64'd47007887360, 64'd13666156, - 64'd1467081088, - 64'd179082544, - 64'd802506014720, 64'd88252309504, 64'd47607111680, 64'd1127799296, - 64'd1363320832, - 64'd196159872, - 64'd838934003712, 64'd57425080320, 64'd47399833600, 64'd2187287808, - 64'd1242587520, - 64'd209838160, - 64'd859940061184, 64'd26651252736, 64'd46415323136, 64'd3177429760, - 64'd1107204736, - 64'd220019792, - 64'd865679441920, - 64'd3558628352, 64'd44694278144, 64'd4085026560, - 64'd959648448, - 64'd226659696, - 64'd856556503040, - 64'd32719437824, 64'd42287857664, 64'd4898542080, - 64'd802507008, - 64'd229765008, - 64'd833210482688, - 64'd60378497024, 64'd39256571904, 64'd5608235008, - 64'd638439104, - 64'd229393904, - 64'd796497477632, - 64'd86121881600, 64'd35669041152, 64'd6206257664, - 64'd470132416, - 64'd225653632, - 64'd747469733888, - 64'd109579927552, 64'd31600689152, 64'd6686722048, - 64'd300262304, - 64'd218697952, - 64'd687352250368, - 64'd130431860736, 64'd27132338176, 64'd7045738496, - 64'd131451952, - 64'd208723776, - 64'd617517285376, - 64'd148409516032, 64'd22348781568, 64'd7281419776, 64'd33766012, - 64'd195967312, - 64'd539457552384, - 64'd163300114432, 64'd17337327616, 64'd7393851392, 64'd192985360, - 64'd180699632, - 64'd454757908480, - 64'd174948057088, 64'd12186329088, 64'd7385038848, 64'd343959488, - 64'd163221824, - 64'd365066518528, - 64'd183255728128, 64'd6983767040, 64'd7258820096, 64'd484631296, - 64'd143859824, - 64'd272065822720, - 64'd188183445504, 64'd1815849472, 64'd7020755456, 64'd613159616, - 64'd122958880, - 64'd177443848192, - 64'd189748363264, - 64'd3234301184, 64'd6677993984, 64'd727941376, - 64'd100877936, - 64'd82866216960, - 64'd188022505472, - 64'd8087886336, 64'd6239116800, 64'd827629760, - 64'd77983912, 64'd10050632704, - 64'd183130112000, - 64'd12671563776, 64'd5713961984, 64'd911148096, - 64'd54645936, 64'd99764699136, - 64'd175244050432, - 64'd16918459392, 64'd5113438208, 64'd977698944, - 64'd31229768, 64'd184831721472, - 64'd164581588992, - 64'd20769056768, 64'd4449323008, 64'd1026768832, - 64'd8092306, 64'd263926185984, - 64'd151399677952, - 64'd24171935744, 64'd3734053376, 64'd1058128640, 64'd14423572, 64'd335859875840, - 64'd135989600256, - 64'd27084365824, 64'd2980513792, 64'd1071829056, 64'd35993872, 64'd399597600768, - 64'd118671261696, - 64'd29472751616, 64'd2201821440, 64'd1068192768, 64'd56317924, 64'd454270091264, - 64'd99787186176, - 64'd31312910336, 64'd1411112448, 64'd1047801408, 64'd75122352, 64'd499183616000, - 64'd79696314368, - 64'd32590198784, 64'd621336384, 64'd1011480128, 64'd92164568, 64'd533826732032, - 64'd58767691776, - 64'd33299482624, - 64'd154943552, 64'd960277760, 64'd107235656, 64'd557873823744, - 64'd37374169088, - 64'd33444954112, - 64'd905737024, 64'd895444608, 64'd120162680, 64'd571185233920, - 64'd15886231552, - 64'd33039812608, - 64'd1619800192, 64'd818407360, 64'd130810440, 64'd573804773376, 64'd5333987328, - 64'd32105801728, - 64'd2286791936, 64'd730742464, 64'd139082496, 64'd565953953792, 64'd25938384896, - 64'd30672625664, - 64'd2897413120, 64'd634146880, 64'd144921664, 64'd548023926784, 64'd45598187520, - 64'd28777254912, - 64'd3443524096, 64'd530409024, 64'd148309872, 64'd520564146176, 64'd64008802304, - 64'd26463137792, - 64'd3918241280, 64'd421377696, 64'd149267344, 64'd484269522944, 64'd80894140416, - 64'd23779321856, - 64'd4316012544, 64'd308932032, 64'd147851344, 64'd439965057024, 64'd96010354688, - 64'd20779517952, - 64'd4632668160, 64'd194951008, 64'd144154208, 64'd388588961792, 64'd109148995584, - 64'd17521113088, - 64'd4865448448, 64'd81284144, 64'd138301056, 64'd331174313984, 64'd120139448320, - 64'd14064135168, - 64'd5013009408, - 64'd30276684, 64'd130446984, 64'd268829605888, 64'd128850771968, - 64'd10470236160, - 64'd5075404800, - 64'd138023792, 64'd120773768, 64'd202718658560, 64'd135192780800, - 64'd6801641472, - 64'd5054048768, - 64'd240358176, 64'd109486384, 64'd134040117248, 64'd139116445696, - 64'd3120139008, - 64'd4951653888, - 64'd335811680, 64'd96809216, 64'd64006848512, 64'd140613697536, 64'd513904608, - 64'd4772154368, - 64'd423066464, 64'd82981984, - 64'd6174270464, 64'd139716444160, 64'd4042478336, - 64'd4520609792, - 64'd500971680, 64'd68255632, - 64'd75322032128, 64'd136495087616, 64'd7410798592, - 64'd4203092992, - 64'd568556992, 64'd52888100, - 64'd142299611136, 64'd131056402432, 64'd10568109056, - 64'd3826567936, - 64'd625043008, 64'd37140108, - 64'd206032109568, 64'd123540840448, 64'd13468387328, - 64'd3398753024, - 64'd669848256, 64'd21271010, - 64'd265522659328, 64'd114119467008, 64'd16070970368, - 64'd2927977984, - 64'd702593088, 64'd5534769, - 64'd319866830848, 64'd102990364672, 64'd18341064704, - 64'd2423034880, - 64'd723099968, - 64'd9823876, - 64'd368265166848, 64'd90374766592, 64'd20250150912, - 64'd1893024640, - 64'd731391104, - 64'd24572992, - 64'd410033782784, 64'd76512894976, 64'd21776293888, - 64'd1347204352, - 64'd727682368, - 64'd38496744, - 64'd444612771840, 64'd61659594752, 64'd22904309760, - 64'd794834368, - 64'd712374656, - 64'd51398352, - 64'd471572283392, 64'd46079827968, 64'd23625850880, - 64'd245030640, - 64'd686042560, - 64'd63102660, - 64'd490616586240, 64'd30044149760, 64'd23939354624, 64'd293377280, - 64'd649420608, - 64'd73458312, - 64'd501585739776, 64'd13824169984, 64'd23849902080, 64'd811979904, - 64'd603387136, - 64'd82339488, - 64'd504454807552, - 64'd2311850496, 64'd23368964096, 64'd1302911104, - 64'd548946496, - 64'd89647192, - 64'd499331366912, - 64'd18103277568, 64'd22514049024, 64'd1758959872, - 64'd487209728, - 64'd95310104, - 64'd486450528256, - 64'd33301121024, 64'd21308276736, 64'd2173667840, - 64'd419373920, - 64'd99284920, - 64'd466168217600, - 64'd47671787520, 64'd19779858432, 64'd2541413888, - 64'd346700928, - 64'd101556320, - 64'd438952525824, - 64'd61000474624, 64'd17961517056, 64'd2857481216, - 64'd270495520, - 64'd102136416, - 64'd405373714432, - 64'd73094193152, 64'd15889840128, 64'd3118109184, - 64'd192083456, - 64'd101063864, - 64'd366092419072, - 64'd83784359936, 64'd13604604928, 64'd3320529664, - 64'd112789768, - 64'd98402488, - 64'd321847099392, - 64'd92928925696, 64'd11148049408, 64'd3462983936, - 64'd33917672, - 64'd94239632, - 64'd273440227328, - 64'd100414029824, 64'd8564135936, 64'd3544725760, 64'd43271628, - 64'd88684120, - 64'd221723901952, - 64'd106155171840, 64'd5897799168, 64'd3566006272, 64'd117577960, - 64'd81863952, - 64'd167584972800, - 64'd110097866752, 64'd3194200576, 64'd3528044544, 64'd187879696, - 64'd73923784, - 64'd111929999360, - 64'd112217784320, 64'd497996768, 64'd3432982528, 64'd253149584, - 64'd65022140, - 64'd55670218752, - 64'd112520486912, - 64'd2147366144, 64'd3283827200, 64'd312468704, - 64'd55328580, 64'd293226432, - 64'd111040561152, - 64'd4700319744, 64'd3084379648, 64'd365038144, - 64'd45020656, 64'd55083495424, - 64'd107840413696, - 64'd7121794560, 64'd2839154688, 64'd410188800, - 64'd34280916, 64'd107861565440, - 64'd103008600064, - 64'd9375787008, 64'd2553288192, 64'd447388512, - 64'd23293848, 64'd157838802944, - 64'd96657784832, - 64'd11429858304, 64'd2232440832, 64'd476246976, - 64'd12242892, 64'd204288475136, - 64'd88922374144, - 64'd13255571456, 64'd1882692224, 64'd496518336, - 64'd1307557, 64'd246555901952, - 64'd79955836928, - 64'd14828847104, 64'd1510434048, 64'd508101280, 64'd9339338, 64'd284067299328, - 64'd69927788544, - 64'd16130240512, 64'd1122258432, 64'd511036928, 64'd19534240, 64'd316337160192, - 64'd59020926976, - 64'd17145144320, 64'd724847744, 64'd505504416, 64'd29125226, 64'd342973808640, - 64'd47427776512, - 64'd17863899136, 64'd324865088, 64'd491814400, 64'd37974108, 64'd363683708928, - 64'd35347369984, - 64'd18281832448, - 64'd71152392, 64'd470400736, 64'd45958284, 64'd378273693696, - 64'd22981933056, - 64'd18399207424, - 64'd456894976, 64'd441810336, 64'd52972284, 64'd386651848704, - 64'd10533573632, - 64'd18221096960, - 64'd826375808, 64'd406691392, 64'd58928988, 64'd388826595328, 64'd1798948096, - 64'd17757192192, - 64'd1174018944, 64'd365780480, 64'd63760556, 64'd384904298496, 64'd13823309824, - 64'd17021529088, - 64'd1494738304, 64'd319888416, 64'd67418992, 64'd375085203456, 64'd25356541952, - 64'd16032155648, - 64'd1784006784, 64'd269885376, 64'd69876376, 64'd359658192896, 64'd36227723264, - 64'd14810752000, - 64'd2037915392, 64'd216685360, 64'd71124832, 64'd338994003968, 64'd46280421376, - 64'd13382192128, - 64'd2253219584, 64'd161230592, 64'd71176072, 64'd313537560576, 64'd55374839808, - 64'd11774067712, - 64'd2427375104, 64'd104475496, 64'd70060744, 64'd283799191552, 64'd63389650944, - 64'd10016183296, - 64'd2558562304, 64'd47371200, 64'd67827424, 64'd250344865792, 64'd70223495168, - 64'd8140022272, - 64'd2645694720, - 64'd9149640, 64'd64541392, 64'd213786034176, 64'd75796103168, - 64'd6178208256, - 64'd2688421120, - 64'd64187332, 64'd60283132, 64'd174768832512, 64'd80049086464, - 64'd4163952384, - 64'd2687111168, - 64'd116888728, 64'd55146664, 64'd133963022336, 64'd82946351104, - 64'd2130511360, - 64'd2642831616, - 64'd166459696, 64'd49237692, 64'd92050849792, 64'd84474118144, - 64'd110653576, - 64'd2557312768, - 64'd212176416, 64'd42671612, 64'd49715904512, 64'd84640620544, 64'd1863850752, - 64'd2432903936, - 64'd253395088, 64'd35571408, 64'd7632287232, 64'd83475464192, 64'd3762712832, - 64'd2272520192, - 64'd289560384, 64'd28065490, - 64'd33545834496, 64'd81028612096, 64'd5557572608, - 64'd2079582848, - 64'd320211968, 64'd20285500, - 64'd73194119168, 64'd77369139200, 64'd7222403072, - 64'd1857950848, - 64'd344989568, 64'd12364129, - 64'd110727217152, 64'd72583659520, 64'd8733871104, - 64'd1611849088, - 64'd363636256, 64'd4432954, - 64'd145607098368, 64'd66774532096, 64'd10071640064, - 64'd1345791744, - 64'd375999936, - 64'd3379635, - 64'd177350426624, 64'd60057858048, 64'd11218626560, - 64'd1064502912, - 64'd382033088, - 64'd10950404, - 64'd205534920704, 64'd52561313792, 64'd12161187840, - 64'd772835904, - 64'd381791072, - 64'd18163128, - 64'd229804539904, 64'd44421840896, 64'd12889261056, - 64'd475692544, - 64'd375428544, - 64'd24910266, - 64'd249873547264, 64'd35783254016, 64'd13396432896, - 64'd177943536, - 64'd363194560, - 64'd31094466, - 64'd265529311232, 64'd26793799680, 64'd13679954944, 64'd115648360, - 64'd345426240, - 64'd36629864, - 64'd276633911296, 64'd17603684352, 64'd13740696576, 64'd400501952, - 64'd322541184, - 64'd41443168, - 64'd283124531200, 64'd8362662400, 64'd13583045632, 64'd672286208, - 64'd295028768, - 64'd45474524, - 64'd285012590592, - 64'd782341184, 64'd13214753792, 64'd926983424, - 64'd263440544, - 64'd48678116, - 64'd282381877248, - 64'd9689481216, 64'd12646726656, 64'd1160945536, - 64'd228379888, - 64'd51022572, - 64'd275385253888, - 64'd18224119808, 64'd11892779008, 64'd1370943232, - 64'd190491040, - 64'd52491072, - 64'd264240807936, - 64'd26260789248, 64'd10969340928, 64'd1554207488, - 64'd150447840, - 64'd53081284, - 64'd249226625024, - 64'd33684951040, 64'd9895136256, 64'd1708462336, - 64'd108942160, - 64'd52805020, - 64'd230675021824, - 64'd40394547200, 64'd8690825216, 64'd1831949184, - 64'd66672452, - 64'd51687692, - 64'd208965959680, - 64'd46301310976, 64'd7378630656, 64'd1923442048, - 64'd24332392, - 64'd49767576, - 64'd184519835648, - 64'd51331833856, 64'd5981947904, 64'd1982254208, 64'd17400088, - 64'd47094876, - 64'd157789880320, - 64'd55428366336, 64'd4524942848, 64'd2008235904, 64'd57873236, - 64'd43730612, - 64'd129254154240, - 64'd58549334016, 64'd3032150016, 64'd2001763840, 64'd96471240, - 64'd39745388, - 64'd99407421440, - 64'd60669616128, 64'd1528072832, 64'd1963721984, 64'd132623208, - 64'd35218024, - 64'd68752859136, - 64'd61780545536, 64'd36796504, 64'd1895475328, 64'd165811136, - 64'd30234082, - 64'd37793939456, - 64'd61889617920, - 64'd1418385152, 64'd1798836224, 64'd195576944, - 64'd24884336, - 64'd7026437632, - 64'd61020004352, - 64'd2815320320, 64'd1676024704, 64'd221528240, - 64'd19263196, 64'd23069216768, - 64'd59209773056, - 64'd4133322240, 64'd1529623168, 64'd243343024, - 64'd13467098, 64'd52035162112, - 64'd56510943232, - 64'd5353462784, 64'd1362526464, 64'd260773104, - 64'd7592925, 64'd79442788352, - 64'd52988293120, - 64'd6458829824, 64'd1177887744, 64'd273646208, - 64'd1736438, 64'd104898797568, - 64'd48718045184, - 64'd7434744832, 64'd979062912, 64'd281866912, 64'd4009222, 64'd128050544640, - 64'd43786350592, - 64'd8268942848, 64'd769551040, 64'd285416224, 64'd9554955, 64'd148590624768, - 64'd38287704064, - 64'd8951707648, 64'd552936192, 64'd284350048, 64'd14817033, 64'd166260588544, - 64'd32323217408, - 64'd9475960832, 64'd332827776, 64'd278796512, 64'd19718296, 64'd180853850112, - 64'd25998870528, - 64'd9837315072, 64'd112802824, 64'd268952064, 64'd24189226, 64'd192217645056, - 64'd19423698944, - 64'd10034070528, - 64'd103650368, 64'd255076688, 64'd28168872, 64'd200254128128, - 64'd12708000768, - 64'd10067181568, - 64'd313185376, 64'd237488272, 64'd31605606, 64'd204920520704, - 64'd5961550848, - 64'd9940171776, - 64'd512647424, 64'd216556032, 64'd34457716, 64'd206228488192, 64'd708124480, - 64'd9659018240, - 64'd699118848, 64'd192693456, 64'd36693844, 64'd204242501632, 64'd7197395456, - 64'd9231992832, - 64'd869959680, 64'd166350592, 64'd38293204, 64'd199077560320, 64'd13408075776, - 64'd8669478912, - 64'd1022842816, 64'd138005968, 64'd39245684, 64'd190896128000, 64'd19248842752, - 64'd7983748096, - 64'd1155783296, 64'd108158320, 64'd39551716, 64'd179904282624, 64'd24636518400, - 64'd7188726272, - 64'd1267161216, 64'd77318152, 64'd39222040, 64'd166347489280, 64'd29497176064, - 64'd6299724288, - 64'd1355739264, 64'd45999272, 64'd38277248, 64'd150505635840, 64'd33767094272, - 64'd5333166592, - 64'd1420672000, 64'd14710599, 64'd36747244, 64'd132687716352, 64'd37393506304, - 64'd4306299904, - 64'd1461510272, - 64'd16051860, 64'd34670516, 64'd113226309632, 64'd40335167488, - 64'd3236899328, - 64'd1478198528, - 64'd45812568, 64'd32093330, 64'd92471631872, 64'd42562719744, - 64'd2142974848, - 64'd1471065856, - 64'd74123520, 64'd29068780, 64'd70785564672, 64'd44058857472, - 64'd1042477568, - 64'd1440811392, - 64'd100570712, 64'd25655798, 64'd48535621632, 64'd44818313216, 64'd46982476, - 64'd1388484224, - 64'd124779864, 64'd21918058, 64'd26089003008, 64'd44847632384, 64'd1108407680, - 64'd1315457664, - 64'd146421424, 64'd17922850, 64'd3806748672, 64'd44164767744, 64'd2125667584, - 64'd1223400064, - 64'd165214688, 64'd13739916, - 64'd17961811968, 64'd42798526464, 64'd3083733504, - 64'd1114240512, - 64'd180931088, 64'd9440287, - 64'd38884319232, 64'd40787836928, 64'd3968889600, - 64'd990132288, - 64'd193396528, 64'd5095112, - 64'd58650222592, 64'd38180864000, 64'd4768918016, - 64'd853412352, - 64'd202492816, 64'd774528, - 64'd76975161344, 64'd35034038272, 64'd5473255936, - 64'd706560576, - 64'd208158176, - 64'd3453433, - 64'd93604839424, 64'd31410925568, 64'd6073121280, - 64'd552156160, - 64'd210386848, - 64'd7523876, - 64'd108318269440, 64'd27381069824, 64'd6561609728, - 64'd392834496, - 64'd209227760, - 64'd11375996, - 64'd120930476032, 64'd23018717184, 64'd6933754880, - 64'd231244032, - 64'd204782480, - 64'd14953949, - 64'd131294502912, 64'd18401529856, 64'd7186563072, - 64'd70003600, - 64'd197202240, - 64'd18207614, - 64'd139302813696, 64'd13609263104, 64'd7319006720, 64'd88338248, - 64'd186684336, - 64'd21093252, - 64'd144888004608, 64'd8722452480, 64'd7331995648, 64'd241342064, - 64'd173467872, - 64'd23574048, - 64'd148022853632, 64'd3821109760, 64'd7228313600, 64'd386713472, - 64'd157828880, - 64'd25620520, - 64'd148719747072, - 64'd1016530176, 64'd7012526592, 64'd522336128, - 64'd140075104, - 64'd27210812, - 64'd147029508096, - 64'd5715210240, 64'd6690865664, 64'd646300800, - 64'd120540240, - 64'd28330850, - 64'd143039594496, - 64'd10203770880, 64'd6271088640, 64'd756930624, - 64'd99578080, - 64'd28974380, - 64'd136871796736, - 64'd14416177152, 64'd5762317312, 64'd852802112, - 64'd77556320, - 64'd29142874, - 64'd128679477248, - 64'd18292439040, 64'd5174857728, 64'd932761088, - 64'd54850424, - 64'd28845310, - 64'd118644285440, - 64'd21779417088, 64'd4520009728, 64'd995934912, - 64'd31837438, - 64'd28097850, - 64'd106972594176, - 64'd24831485952, 64'd3809860352, 64'd1041738880, - 64'd8889991, - 64'd26923408, - 64'd93891592192, - 64'd27411083264, 64'd3057072896, 64'd1069878528, 64'd13629545, - 64'd25351112, - 64'd79645155328, - 64'd29489094656, 64'd2274671616, 64'd1080347136, 64'd35374540, - 64'd23415698, - 64'd64489545728, - 64'd31045109760, 64'd1475826304, 64'd1073418880, 64'd56019228, - 64'd21156812, - 64'd48689025024, - 64'd32067528704, 64'd673638400, 64'd1049637120, 64'd75263368, - 64'd18618256, - 64'd32511469568, - 64'd32553523200, - 64'd119064600, 64'd1009799232, 64'd92836392, - 64'd15847203, - 64'd16223992832, - 64'd32508864512, - 64'd889926592, 64'd954937920, 64'd108500936, - 64'd12893350, - 64'd88746856, - 64'd31947616256, - 64'd1627247104, 64'd886298624, 64'd122055824, - 64'd9808074, 64'd15641138176, - 64'd30891702272, - 64'd2320150784, 64'd805314432, 64'd133338360, - 64'd6643568, 64'd30725345280, - 64'd29370359808, - 64'd2958740480, 64'd713579008, 64'd142225952, - 64'd3452002, 64'd44939878400, - 64'd27419498496, - 64'd3534228480, 64'd612817024, 64'd148637040, - 64'd284680, 64'd58080198656, - 64'd25080952832, - 64'd4039049984, 64'd504853440, 64'd152531456, 64'd2808740, 64'd69964013568, - 64'd22401675264, - 64'd4466952192, 64'd391582240, 64'd153909936, 64'd5781004, 64'd80433602560, - 64'd19432865792, - 64'd4813060608, 64'd274934528, 64'd152813168, 64'd8587947, 64'd89357697024, - 64'd16229040128, - 64'd5073922560, 64'd156846864, 64'd149320128, 64'd11189123, 64'd96632946688, - 64'd12847086592, - 64'd5247527424, 64'd39230476, 64'd143545872, 64'd13548353, 64'd102184812544, - 64'd9345304576, - 64'd5333300736, - 64'd76058528, 64'd135638800, 64'd15634194, 64'd105968074752, - 64'd5782438912, - 64'd5332078080, - 64'd187247280, 64'd125777552, 64'd17420324, 64'd107966783488, - 64'd2216733952, - 64'd5246058496, - 64'd292672224, 64'd114167280, 64'd18885832, 64'd108193816576, 64'd1294978432, - 64'd5078732800, - 64'd390802848, 64'd101035864, 64'd20015412, 64'd106689912832, 64'd4698147328, - 64'd4834797056, - 64'd480262688, 64'd86629656, 64'd20799476, 64'd103522353152, 64'd7941314048, - 64'd4520049152, - 64'd559847360, 64'd71209128, 64'd21234158, 64'd98783232000, 64'd10976852992, - 64'd4141266432, - 64'd628539328, 64'd55044372, 64'd21321234, 64'd92587327488, 64'd13761633280, - 64'd3706075648, - 64'd685519616, 64'd38410596, 64'd21067960, 64'd85069766656, 64'd16257591296, - 64'd3222810112, - 64'd730175616, 64'd21583592, 64'd20486812, 64'd76383322112, 64'd18432212992, - 64'd2700358656, - 64'd762106048, 64'd4835369, 64'd19595166, 64'd66695573504, 64'd20258908160, - 64'd2148011520, - 64'd781121600, - 64'd11570094, 64'd18414896, 64'd56185835520, 64'd21717288960, - 64'd1575302784, - 64'd787243072, - 64'd27380832, 64'd16971916, 64'd45042040832, 64'd22793334784, - 64'd991851136, - 64'd780695552, - 64'd42360600, 64'd15295670, 64'd33457522688, 64'd23479463936, - 64'd407206720, - 64'd761899904, - 64'd56292244, 64'd13418574, 64'd21627799552, 64'd23774482432, 64'd169300192, - 64'd731461184, - 64'd68980656, 64'd11375428, 64'd9747416064, 64'd23683454976, 64'd728701632, - 64'd690154240, - 64'd80255344, 64'd9202805, - 64'd1993129344, 64'd23217463296, 64'd1262525568, - 64'd638907456, - 64'd89972536, 64'd6938424, - 64'd13410318336, 64'd22393276416, 64'd1762918144, - 64'd578783936, - 64'd98016768, 64'd4620524, - 64'd24330354688, 64'd21232945152, 64'd2222753536, - 64'd510961472, - 64'd104302040, 64'd2287246, - 64'd34591690752, 64'd19763324928, 64'd2635728128, - 64'd436710720, - 64'd108772432, - 64'd23980, - 64'd44047294464, 64'd18015514624, 64'd2996441856, - 64'd357372896, - 64'd111402280, - 64'd2276999, - 64'd52566618112, 64'd16024272896, 64'd3300460032, - 64'd274336512, - 64'd112195776, - 64'd4437484, - 64'd60037275648, 64'd13827361792, 64'd3544360448, - 64'd189014320, - 64'd111186200, - 64'd6473431, - 64'd66366373888, 64'd11464875008, 64'd3725762560, - 64'd102820136, - 64'd108434648, - 64'd8355611, - 64'd71481499648, 64'd8978542592, 64'd3843339264, - 64'd17146324, - 64'd104028384, - 64'd10057966, - 64'd75331379200, 64'd6411025408, 64'd3896812032, 64'd66657732, - 64'd98078776, - 64'd11557943, - 64'd77886144512, 64'd3805214208, 64'd3886928128, 64'd147306064, - 64'd90718944, - 64'd12836766, - 64'd79137292288, 64'd1203540608, 64'd3815425280, 64'd223594944, - 64'd82101112, - 64'd13879640, - 64'd79097274368, - 64'd1352686720, 64'd3684976896, 64'd294420000, - 64'd72393696, - 64'd14675887, - 64'd77798785024, - 64'd3823910656, 64'd3499128064, 64'd358791296, - 64'd61778220, - 64'd15219014, - 64'd75293745152, - 64'd6172911616, 64'd3262216448, 64'd415846208, - 64'd50446116, - 64'd15506713, - 64'd71651991552, - 64'd8365341184, 64'd2979283968, 64'd464859936, - 64'd38595436, - 64'd15540788, - 64'd66959687680, - 64'd10370196480, 64'd2655979008, 64'd505253664, - 64'd26427528, - 64'd15327032, - 64'd61317615616, - 64'd12160233472, 64'd2298451200, 64'd536600032, - 64'd14143770, - 64'd14875031, - 64'd54839140352, - 64'd13712301056, 64'd1913241984, 64'd558626304, - 64'd1942347, - 64'd14197915, - 64'd47648133120, - 64'd15007612928, 64'd1507169536, 64'd571214592, 64'd9984802, - 64'd13312069, - 64'd39876722688, - 64'd16031933440, 64'd1087214208, 64'd574400256, 64'd21454888, - 64'd12236782, - 64'd31662987264, - 64'd16775695360, 64'd660403712, 64'd568367104, 64'd32296946, - 64'd10993875, - 64'd23148623872, - 64'd17234030592, 64'd233699392, 64'd553441088, 64'd42354264, - 64'd9607290, - 64'd14476587008, - 64'd17406736384, - 64'd186112288, 64'd530081408, 64'd51486508, - 64'd8102654, - 64'd5788791296, - 64'd17298159616, - 64'd592523456, 64'd498869920, 64'd59571556, - 64'd6506830, 64'd2776121088, - 64'd16917010432, - 64'd979401536, 64'd460498944, 64'd66506984, - 64'd4847465, 64'd11084907520, - 64'd16276123648, - 64'd1341077248, 64'd415757280, 64'd72211192, - 64'd3152522, 64'd19011708928, - 64'd15392145408, - 64'd1672423168, 64'd365515520, 64'd76624208, - 64'd1449835, 64'd26439870464, - 64'd14285174784, - 64'd1968922496, 64'd310709952, 64'd79708064, 64'd233334, 64'd33263562752, - 64'd12978362368, - 64'd2226724608, 64'd252326112, 64'd81446888, 64'd1870714, 64'd39389204480, - 64'd11497459712, - 64'd2442690560, 64'd191381936, 64'd81846584, 64'd3437414, 64'd44736643072, - 64'd9870348288, - 64'd2614424576, 64'd128910704, 64'd80934216, 64'd4910289};
endpackage
`endif
