`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam N = 4;
	localparam M = 4;
	localparam real Lfr[0:3] = {0.98044646, 0.98044646, 0.9601575, 0.9601575};
	localparam real Lfi[0:3] = {0.07935079, -0.07935079, 0.03143782, -0.03143782};
	localparam real Lbr[0:3] = {0.98044646, 0.98044646, 0.9601575, 0.9601575};
	localparam real Lbi[0:3] = {0.07935079, -0.07935079, 0.03143782, -0.03143782};
	localparam real Wfr[0:3] = {0.000101395075, 0.000101395075, 2.9913577e-05, 2.9913577e-05};
	localparam real Wfi[0:3] = {5.1355123e-06, -5.1355123e-06, 5.8664347e-05, -5.8664347e-05};
	localparam real Wbr[0:3] = {-0.000101395075, -0.000101395075, -2.9913577e-05, -2.9913577e-05};
	localparam real Wbi[0:3] = {-5.1355123e-06, 5.1355123e-06, -5.8664347e-05, 5.8664347e-05};
	localparam real Ffr[0:3][0:79] = '{
		'{40.21009, 6.34191, -1.2044557, 0.02154542, 43.19078, 5.5783777, -1.212442, 0.032587305, 45.786346, 4.8023486, -1.2120714, 0.04305347, 47.99194, 4.01941, -1.2036176, 0.052892692, 49.805477, 3.2350156, -1.1873991, 0.06205958, 51.22756, 2.4544513, -1.163776, 0.070514716, 52.261383, 1.6828065, -1.1331463, 0.0782247, 52.912636, 0.92494524, -1.0959415, 0.085162215, 53.18937, 0.18548255, -1.0526237, 0.09130597, 53.101883, -0.53123957, -1.0036802, 0.09664067, 52.662575, -1.2211715, -0.9496205, 0.10115692, 51.88578, -1.8805742, -0.8909713, 0.104851104, 50.78764, -2.5060334, -0.82827336, 0.1077252, 49.385906, -3.094473, -0.7620766, 0.109786615, 47.699783, -3.6431625, -0.6929367, 0.11104793, 45.749756, -4.149727, -0.62141085, 0.11152666, 43.557407, -4.6121483, -0.5480541, 0.111245, 41.14524, -5.028771, -0.47341576, 0.11022947, 38.536488, -5.398296, -0.39803594, 0.108510666, 35.75495, -5.719784, -0.3224421, 0.10612287},
		'{40.21009, 6.34191, -1.2044557, 0.02154542, 43.19078, 5.5783777, -1.212442, 0.032587305, 45.786346, 4.8023486, -1.2120714, 0.04305347, 47.99194, 4.01941, -1.2036176, 0.052892692, 49.805477, 3.2350156, -1.1873991, 0.06205958, 51.22756, 2.4544513, -1.163776, 0.070514716, 52.261383, 1.6828065, -1.1331463, 0.0782247, 52.912636, 0.92494524, -1.0959415, 0.085162215, 53.18937, 0.18548255, -1.0526237, 0.09130597, 53.101883, -0.53123957, -1.0036802, 0.09664067, 52.662575, -1.2211715, -0.9496205, 0.10115692, 51.88578, -1.8805742, -0.8909713, 0.104851104, 50.78764, -2.5060334, -0.82827336, 0.1077252, 49.385906, -3.094473, -0.7620766, 0.109786615, 47.699783, -3.6431625, -0.6929367, 0.11104793, 45.749756, -4.149727, -0.62141085, 0.11152666, 43.557407, -4.6121483, -0.5480541, 0.111245, 41.14524, -5.028771, -0.47341576, 0.11022947, 38.536488, -5.398296, -0.39803594, 0.108510666, 35.75495, -5.719784, -0.3224421, 0.10612287},
		'{39.456413, 6.232743, -1.1224245, 0.2605331, 42.39817, 5.5410104, -1.0205656, 0.2445576, 45.003883, 4.888345, -0.9239323, 0.22918406, 47.29275, 4.273414, -0.83237046, 0.21440563, 49.283314, 3.6948936, -0.7457249, 0.2002145, 50.993443, 3.1514647, -0.6638397, 0.18660194, 52.440357, 2.641822, -0.58655876, 0.17355837, 53.64063, 2.1646726, -0.513726, 0.16107355, 54.610184, 1.7187403, -0.44518608, 0.14913653, 55.36431, 1.3027663, -0.38078454, 0.13773583, 55.917686, 0.9155122, -0.32036814, 0.12685946, 56.28436, 0.55576074, -0.2637852, 0.11649499, 56.477787, 0.22231795, -0.2108859, 0.106629655, 56.510822, -0.08598599, -0.16152242, 0.09725038, 56.395752, -0.37029538, -0.115549274, 0.08834383, 56.144295, -0.6317281, -0.07282345, 0.07989651, 55.767612, -0.8713748, -0.033204608, 0.071894765, 55.27633, -1.090298, 0.0034447827, 0.06432484, 54.680553, -1.289532, 0.037259296, 0.057172943, 53.989872, -1.4700816, 0.06837043, 0.050425258},
		'{39.456413, 6.232743, -1.1224245, 0.2605331, 42.39817, 5.5410104, -1.0205656, 0.2445576, 45.003883, 4.888345, -0.9239323, 0.22918406, 47.29275, 4.273414, -0.83237046, 0.21440563, 49.283314, 3.6948936, -0.7457249, 0.2002145, 50.993443, 3.1514647, -0.6638397, 0.18660194, 52.440357, 2.641822, -0.58655876, 0.17355837, 53.64063, 2.1646726, -0.513726, 0.16107355, 54.610184, 1.7187403, -0.44518608, 0.14913653, 55.36431, 1.3027663, -0.38078454, 0.13773583, 55.917686, 0.9155122, -0.32036814, 0.12685946, 56.28436, 0.55576074, -0.2637852, 0.11649499, 56.477787, 0.22231795, -0.2108859, 0.106629655, 56.510822, -0.08598599, -0.16152242, 0.09725038, 56.395752, -0.37029538, -0.115549274, 0.08834383, 56.144295, -0.6317281, -0.07282345, 0.07989651, 55.767612, -0.8713748, -0.033204608, 0.071894765, 55.27633, -1.090298, 0.0034447827, 0.06432484, 54.680553, -1.289532, 0.037259296, 0.057172943, 53.989872, -1.4700816, 0.06837043, 0.050425258}};
	localparam real Ffi[0:3][0:79] = '{
		'{-47.47199, 8.059468, 0.3974449, -0.14446199, -43.35304, 8.405112, 0.2940989, -0.1399276, -39.078114, 8.683412, 0.19214001, -0.13460569, -34.680813, 8.8946905, 0.09220417, -0.12855735, -30.194483, 9.039711, -0.00510676, -0.12184652, -25.65197, 9.119654, -0.099227965, -0.11453951, -21.085436, 9.136095, -0.18963425, -0.10670446, -16.526157, 9.090983, -0.27584228, -0.09841082, -12.004354, 8.986618, -0.35741243, -0.08972885, -7.5490074, 8.825616, -0.43395028, -0.080729134, -3.187721, 8.610889, -0.5051078, -0.07148208, 1.0534272, 8.345615, -0.57058436, -0.06205747, 5.150007, 8.033204, -0.63012666, -0.052524004, 9.079346, 7.6772704, -0.6835296, -0.042948894, 12.820622, 7.281604, -0.7306356, -0.033397436, 16.35495, 6.850135, -0.7713341, -0.023932658, 19.665432, 6.386906, -0.80556124, -0.01461496, 22.737219, 5.896042, -0.8332982, -0.005501807, 25.557533, 5.3817167, -0.8545702, 0.0033525687, 28.115692, 4.848126, -0.8694448, 0.011897421},
		'{47.47199, -8.059468, -0.3974449, 0.14446199, 43.35304, -8.405112, -0.2940989, 0.1399276, 39.078114, -8.683412, -0.19214001, 0.13460569, 34.680813, -8.8946905, -0.09220417, 0.12855735, 30.194483, -9.039711, 0.00510676, 0.12184652, 25.65197, -9.119654, 0.099227965, 0.11453951, 21.085436, -9.136095, 0.18963425, 0.10670446, 16.526157, -9.090983, 0.27584228, 0.09841082, 12.004354, -8.986618, 0.35741243, 0.08972885, 7.5490074, -8.825616, 0.43395028, 0.080729134, 3.187721, -8.610889, 0.5051078, 0.07148208, -1.0534272, -8.345615, 0.57058436, 0.06205747, -5.150007, -8.033204, 0.63012666, 0.052524004, -9.079346, -7.6772704, 0.6835296, 0.042948894, -12.820622, -7.281604, 0.7306356, 0.033397436, -16.35495, -6.850135, 0.7713341, 0.023932658, -19.665432, -6.386906, 0.80556124, 0.01461496, -22.737219, -5.896042, 0.8332982, 0.005501807, -25.557533, -5.3817167, 0.8545702, -0.0033525687, -28.115692, -4.848126, 0.8694448, -0.011897421},
		'{-143.5786, 14.104169, -1.8175136, 0.17797658, -136.61765, 13.738168, -1.780386, 0.17907615, -129.84155, 13.365002, -1.7415353, 0.17962967, -123.253525, 12.986186, -1.7011946, 0.17967781, -116.85602, 12.603131, -1.6595827, 0.17925946, -110.65082, 12.217151, -1.6169049, 0.17841162, -104.6391, 11.829464, -1.573353, 0.17716962, -98.8214, 11.441202, -1.5291069, 0.17556705, -93.19777, 11.053409, -1.4843339, 0.17363581, -87.767715, 10.667047, -1.43919, 0.17140627, -82.5303, 10.283002, -1.3938202, 0.16890712, -77.48415, 9.902083, -1.3483586, 0.16616563, -72.62754, 9.525031, -1.3029295, 0.16320753, -67.958336, 9.152519, -1.2576473, 0.16005714, -63.474133, 8.785157, -1.2126174, 0.1567374, -59.172207, 8.423493, -1.1679363, 0.15326993, -55.049583, 8.068021, -1.1236923, 0.14967506, -51.103058, 7.7191763, -1.0799655, 0.14597185, -47.32922, 7.377349, -1.0368286, 0.1421782, -43.72447, 7.0428767, -0.9943475, 0.13831086},
		'{143.5786, -14.104169, 1.8175136, -0.17797658, 136.61765, -13.738168, 1.780386, -0.17907615, 129.84155, -13.365002, 1.7415353, -0.17962967, 123.253525, -12.986186, 1.7011946, -0.17967781, 116.85602, -12.603131, 1.6595827, -0.17925946, 110.65082, -12.217151, 1.6169049, -0.17841162, 104.6391, -11.829464, 1.573353, -0.17716962, 98.8214, -11.441202, 1.5291069, -0.17556705, 93.19777, -11.053409, 1.4843339, -0.17363581, 87.767715, -10.667047, 1.43919, -0.17140627, 82.5303, -10.283002, 1.3938202, -0.16890712, 77.48415, -9.902083, 1.3483586, -0.16616563, 72.62754, -9.525031, 1.3029295, -0.16320753, 67.958336, -9.152519, 1.2576473, -0.16005714, 63.474133, -8.785157, 1.2126174, -0.1567374, 59.172207, -8.423493, 1.1679363, -0.15326993, 55.049583, -8.068021, 1.1236923, -0.14967506, 51.103058, -7.7191763, 1.0799655, -0.14597185, 47.32922, -7.377349, 1.0368286, -0.1421782, 43.72447, -7.0428767, 0.9943475, -0.13831086}};
	localparam real Fbr[0:3][0:79] = '{
		'{-40.21009, 6.34191, 1.2044557, 0.02154542, -43.19078, 5.5783777, 1.212442, 0.032587305, -45.786346, 4.8023486, 1.2120714, 0.04305347, -47.99194, 4.01941, 1.2036176, 0.052892692, -49.805477, 3.2350156, 1.1873991, 0.06205958, -51.22756, 2.4544513, 1.163776, 0.070514716, -52.261383, 1.6828065, 1.1331463, 0.0782247, -52.912636, 0.92494524, 1.0959415, 0.085162215, -53.18937, 0.18548255, 1.0526237, 0.09130597, -53.101883, -0.53123957, 1.0036802, 0.09664067, -52.662575, -1.2211715, 0.9496205, 0.10115692, -51.88578, -1.8805742, 0.8909713, 0.104851104, -50.78764, -2.5060334, 0.82827336, 0.1077252, -49.385906, -3.094473, 0.7620766, 0.109786615, -47.699783, -3.6431625, 0.6929367, 0.11104793, -45.749756, -4.149727, 0.62141085, 0.11152666, -43.557407, -4.6121483, 0.5480541, 0.111245, -41.14524, -5.028771, 0.47341576, 0.11022947, -38.536488, -5.398296, 0.39803594, 0.108510666, -35.75495, -5.719784, 0.3224421, 0.10612287},
		'{-40.21009, 6.34191, 1.2044557, 0.02154542, -43.19078, 5.5783777, 1.212442, 0.032587305, -45.786346, 4.8023486, 1.2120714, 0.04305347, -47.99194, 4.01941, 1.2036176, 0.052892692, -49.805477, 3.2350156, 1.1873991, 0.06205958, -51.22756, 2.4544513, 1.163776, 0.070514716, -52.261383, 1.6828065, 1.1331463, 0.0782247, -52.912636, 0.92494524, 1.0959415, 0.085162215, -53.18937, 0.18548255, 1.0526237, 0.09130597, -53.101883, -0.53123957, 1.0036802, 0.09664067, -52.662575, -1.2211715, 0.9496205, 0.10115692, -51.88578, -1.8805742, 0.8909713, 0.104851104, -50.78764, -2.5060334, 0.82827336, 0.1077252, -49.385906, -3.094473, 0.7620766, 0.109786615, -47.699783, -3.6431625, 0.6929367, 0.11104793, -45.749756, -4.149727, 0.62141085, 0.11152666, -43.557407, -4.6121483, 0.5480541, 0.111245, -41.14524, -5.028771, 0.47341576, 0.11022947, -38.536488, -5.398296, 0.39803594, 0.108510666, -35.75495, -5.719784, 0.3224421, 0.10612287},
		'{-39.456413, 6.232743, 1.1224245, 0.2605331, -42.39817, 5.5410104, 1.0205656, 0.2445576, -45.003883, 4.888345, 0.9239323, 0.22918406, -47.29275, 4.273414, 0.83237046, 0.21440563, -49.283314, 3.6948936, 0.7457249, 0.2002145, -50.993443, 3.1514647, 0.6638397, 0.18660194, -52.440357, 2.641822, 0.58655876, 0.17355837, -53.64063, 2.1646726, 0.513726, 0.16107355, -54.610184, 1.7187403, 0.44518608, 0.14913653, -55.36431, 1.3027663, 0.38078454, 0.13773583, -55.917686, 0.9155122, 0.32036814, 0.12685946, -56.28436, 0.55576074, 0.2637852, 0.11649499, -56.477787, 0.22231795, 0.2108859, 0.106629655, -56.510822, -0.08598599, 0.16152242, 0.09725038, -56.395752, -0.37029538, 0.115549274, 0.08834383, -56.144295, -0.6317281, 0.07282345, 0.07989651, -55.767612, -0.8713748, 0.033204608, 0.071894765, -55.27633, -1.090298, -0.0034447827, 0.06432484, -54.680553, -1.289532, -0.037259296, 0.057172943, -53.989872, -1.4700816, -0.06837043, 0.050425258},
		'{-39.456413, 6.232743, 1.1224245, 0.2605331, -42.39817, 5.5410104, 1.0205656, 0.2445576, -45.003883, 4.888345, 0.9239323, 0.22918406, -47.29275, 4.273414, 0.83237046, 0.21440563, -49.283314, 3.6948936, 0.7457249, 0.2002145, -50.993443, 3.1514647, 0.6638397, 0.18660194, -52.440357, 2.641822, 0.58655876, 0.17355837, -53.64063, 2.1646726, 0.513726, 0.16107355, -54.610184, 1.7187403, 0.44518608, 0.14913653, -55.36431, 1.3027663, 0.38078454, 0.13773583, -55.917686, 0.9155122, 0.32036814, 0.12685946, -56.28436, 0.55576074, 0.2637852, 0.11649499, -56.477787, 0.22231795, 0.2108859, 0.106629655, -56.510822, -0.08598599, 0.16152242, 0.09725038, -56.395752, -0.37029538, 0.115549274, 0.08834383, -56.144295, -0.6317281, 0.07282345, 0.07989651, -55.767612, -0.8713748, 0.033204608, 0.071894765, -55.27633, -1.090298, -0.0034447827, 0.06432484, -54.680553, -1.289532, -0.037259296, 0.057172943, -53.989872, -1.4700816, -0.06837043, 0.050425258}};
	localparam real Fbi[0:3][0:79] = '{
		'{47.47199, 8.059468, -0.3974449, -0.14446199, 43.35304, 8.405112, -0.2940989, -0.1399276, 39.078114, 8.683412, -0.19214001, -0.13460569, 34.680813, 8.8946905, -0.09220417, -0.12855735, 30.194483, 9.039711, 0.00510676, -0.12184652, 25.65197, 9.119654, 0.099227965, -0.11453951, 21.085436, 9.136095, 0.18963425, -0.10670446, 16.526157, 9.090983, 0.27584228, -0.09841082, 12.004354, 8.986618, 0.35741243, -0.08972885, 7.5490074, 8.825616, 0.43395028, -0.080729134, 3.187721, 8.610889, 0.5051078, -0.07148208, -1.0534272, 8.345615, 0.57058436, -0.06205747, -5.150007, 8.033204, 0.63012666, -0.052524004, -9.079346, 7.6772704, 0.6835296, -0.042948894, -12.820622, 7.281604, 0.7306356, -0.033397436, -16.35495, 6.850135, 0.7713341, -0.023932658, -19.665432, 6.386906, 0.80556124, -0.01461496, -22.737219, 5.896042, 0.8332982, -0.005501807, -25.557533, 5.3817167, 0.8545702, 0.0033525687, -28.115692, 4.848126, 0.8694448, 0.011897421},
		'{-47.47199, -8.059468, 0.3974449, 0.14446199, -43.35304, -8.405112, 0.2940989, 0.1399276, -39.078114, -8.683412, 0.19214001, 0.13460569, -34.680813, -8.8946905, 0.09220417, 0.12855735, -30.194483, -9.039711, -0.00510676, 0.12184652, -25.65197, -9.119654, -0.099227965, 0.11453951, -21.085436, -9.136095, -0.18963425, 0.10670446, -16.526157, -9.090983, -0.27584228, 0.09841082, -12.004354, -8.986618, -0.35741243, 0.08972885, -7.5490074, -8.825616, -0.43395028, 0.080729134, -3.187721, -8.610889, -0.5051078, 0.07148208, 1.0534272, -8.345615, -0.57058436, 0.06205747, 5.150007, -8.033204, -0.63012666, 0.052524004, 9.079346, -7.6772704, -0.6835296, 0.042948894, 12.820622, -7.281604, -0.7306356, 0.033397436, 16.35495, -6.850135, -0.7713341, 0.023932658, 19.665432, -6.386906, -0.80556124, 0.01461496, 22.737219, -5.896042, -0.8332982, 0.005501807, 25.557533, -5.3817167, -0.8545702, -0.0033525687, 28.115692, -4.848126, -0.8694448, -0.011897421},
		'{143.5786, 14.104169, 1.8175136, 0.17797658, 136.61765, 13.738168, 1.780386, 0.17907615, 129.84155, 13.365002, 1.7415353, 0.17962967, 123.253525, 12.986186, 1.7011946, 0.17967781, 116.85602, 12.603131, 1.6595827, 0.17925946, 110.65082, 12.217151, 1.6169049, 0.17841162, 104.6391, 11.829464, 1.573353, 0.17716962, 98.8214, 11.441202, 1.5291069, 0.17556705, 93.19777, 11.053409, 1.4843339, 0.17363581, 87.767715, 10.667047, 1.43919, 0.17140627, 82.5303, 10.283002, 1.3938202, 0.16890712, 77.48415, 9.902083, 1.3483586, 0.16616563, 72.62754, 9.525031, 1.3029295, 0.16320753, 67.958336, 9.152519, 1.2576473, 0.16005714, 63.474133, 8.785157, 1.2126174, 0.1567374, 59.172207, 8.423493, 1.1679363, 0.15326993, 55.049583, 8.068021, 1.1236923, 0.14967506, 51.103058, 7.7191763, 1.0799655, 0.14597185, 47.32922, 7.377349, 1.0368286, 0.1421782, 43.72447, 7.0428767, 0.9943475, 0.13831086},
		'{-143.5786, -14.104169, -1.8175136, -0.17797658, -136.61765, -13.738168, -1.780386, -0.17907615, -129.84155, -13.365002, -1.7415353, -0.17962967, -123.253525, -12.986186, -1.7011946, -0.17967781, -116.85602, -12.603131, -1.6595827, -0.17925946, -110.65082, -12.217151, -1.6169049, -0.17841162, -104.6391, -11.829464, -1.573353, -0.17716962, -98.8214, -11.441202, -1.5291069, -0.17556705, -93.19777, -11.053409, -1.4843339, -0.17363581, -87.767715, -10.667047, -1.43919, -0.17140627, -82.5303, -10.283002, -1.3938202, -0.16890712, -77.48415, -9.902083, -1.3483586, -0.16616563, -72.62754, -9.525031, -1.3029295, -0.16320753, -67.958336, -9.152519, -1.2576473, -0.16005714, -63.474133, -8.785157, -1.2126174, -0.1567374, -59.172207, -8.423493, -1.1679363, -0.15326993, -55.049583, -8.068021, -1.1236923, -0.14967506, -51.103058, -7.7191763, -1.0799655, -0.14597185, -47.32922, -7.377349, -1.0368286, -0.1421782, -43.72447, -7.0428767, -0.9943475, -0.13831086}};
	localparam real hf[0:1199] = {0.027848251, -7.863854e-05, -0.000102238904, 5.581651e-07, 0.027769677, -0.00023546736, -0.000101059166, 1.6659997e-06, 0.027612986, -0.000390961, -9.87138e-05, 2.7490748e-06, 0.027379066, -0.0005442468, -9.5228235e-05, 3.7924478e-06, 0.027069231, -0.0006944717, -9.0638314e-05, 4.7825465e-06, 0.026685225, -0.00084080873, -8.498945e-05, 5.7071875e-06, 0.026229188, -0.0009824634, -7.833585e-05, 6.5555873e-06, 0.025703654, -0.001118679, -7.073963e-05, 7.3183596e-06, 0.02511152, -0.0012487425, -6.227e-05, 7.98751e-06, 0.024456035, -0.0013719881, -5.300233e-05, 8.556417e-06, 0.023740761, -0.0014878028, -4.301732e-05, 9.01981e-06, 0.022969553, -0.0015956288, -3.240009e-05, 9.373733e-06, 0.022146536, -0.0016949669, -2.1239324e-05, 9.615509e-06, 0.021276066, -0.0017853795, -9.626397e-06, 9.743692e-06, 0.0203627, -0.0018664917, 2.3454697e-06, 9.758017e-06, 0.019411169, -0.0019379936, 1.4582022e-05, 9.659341e-06, 0.018426342, -0.0019996406, 2.698878e-05, 9.449581e-06, 0.017413195, -0.0020512538, 3.9471804e-05, 9.131647e-06, 0.016376775, -0.0020927207, 5.193842e-05, 8.709373e-06, 0.01532217, -0.0021239934, 6.429791e-05, 8.187441e-06, 0.014254476, -0.0021450883, 7.646218e-05, 7.5713097e-06, 0.013178764, -0.0021560842, 8.834636e-05, 6.8671284e-06, 0.01210005, -0.0021571212, 9.9869336e-05, 6.0816633e-06, 0.011023269, -0.0021483973, 0.00011095432, 5.2222153e-06, 0.009953238, -0.0021301666, 0.000121529265, 4.296539e-06, 0.008894636, -0.0021027357, 0.00013152728, 3.3127621e-06, 0.007851977, -0.0020664614, 0.000140887, 2.2793056e-06, 0.006829583, -0.0020217458, 0.00014955288, 1.2048044e-06, 0.005831566, -0.0019690336, 0.00015747549, 9.803153e-08, 0.004861804, -0.0019088082, 0.0001646116, -1.0321777e-06, 0.0039239265, -0.001841587, 0.00017092444, -2.176997e-06, 0.0030212952, -0.0017679174, 0.00017638376, -3.3276792e-06, 0.0021569917, -0.0016883726, 0.00018096587, -4.4756216e-06, 0.0013338061, -0.0016035473, 0.00018465356, -5.6124286e-06, 0.0005542263, -0.001514053, 0.0001874362, -6.7299707e-06, -0.00017956895, -0.0014205141, 0.00018930952, -7.820437e-06, -0.00086571515, -0.0013235628, 0.00019027547, -8.876385e-06, -0.0015026652, -0.0012238359, 0.00019034215, -9.890792e-06, -0.0020891905, -0.0011219693, 0.00018952347, -1.0857087e-05, -0.0026243792, -0.001018595, 0.00018783894, -1.176919e-05, -0.0031076341, -0.00091433653, 0.00018531342, -1.26215455e-05, -0.0035386665, -0.0008098057, 0.00018197673, -1.3409146e-05, -0.00391749, -0.00070559845, 0.0001778634, -1.4127555e-05, -0.0042444114, -0.0006022919, 0.00017301223, -1.477292e-05, -0.0045200214, -0.00050044095, 0.00016746596, -1.5341988e-05, -0.0047451803, -0.00040057558, 0.00016127084, -1.5832109e-05, -0.0049210084, -0.0003031979, 0.00015447625, -1.6241243e-05, -0.0050488687, -0.00020878005, 0.00014713424, -1.6567954e-05, -0.0051303525, -0.00011776187, 0.00013929917, -1.6811402e-05, -0.0051672626, -3.0549036e-05, 0.0001310272, -1.6971335e-05, -0.0051615955, 5.2488434e-05, 0.00012237595, -1.7048078e-05, -0.0051155235, 0.00013101756, 0.000113403985, -1.7042508e-05, -0.005031377, 0.00020474338, 0.00010417048, -1.6956043e-05, -0.0049116225, 0.00027340974, 9.473475e-05, -1.6790598e-05, -0.0047588455, 0.00033679965, 8.515589e-05, -1.6548585e-05, -0.0045757308, 0.00039473572, 7.549234e-05, -1.6232862e-05, -0.0043650414, 0.00044707974, 6.580157e-05, -1.5846703e-05, -0.0041295993, 0.0004937327, 5.6139706e-05, -1.539378e-05, -0.0038722672, 0.000534634, 4.656119e-05, -1.4878104e-05, -0.0035959282, 0.0005697608, 3.711847e-05, -1.4304009e-05, -0.003303467, 0.00059912674, 2.7861719e-05, -1.3676101e-05, -0.002997754, 0.00062278105, 1.8838567e-05, -1.2999224e-05, -0.002681625, 0.0006408069, 1.0093863e-05, -1.2278419e-05, -0.002357867, 0.0006533199, 1.6694551e-06, -1.1518884e-05, -0.0020292008, 0.00066046615, -6.395991e-06, -1.072594e-05, -0.0016982675, 0.0006624206, -1.4067155e-05, -9.904985e-06, -0.0013676136, 0.0006593847, -2.1312191e-05, -9.0614585e-06, -0.0010396786, 0.0006515847, -2.8102844e-05, -8.200804e-06, -0.0007167833, 0.00063926884, -3.441452e-05, -7.3284336e-06, -0.00040111947, 0.0006227055, -4.0226332e-05, -6.4496917e-06, -9.4740004e-05, 0.00060218055, -4.5521145e-05, -5.5698206e-06, 0.00020044901, 0.0005779951, -5.028556e-05, -4.6939313e-06, 0.0004826953, 0.0005504629, -5.4509896e-05, -3.826971e-06, 0.0007504061, 0.00051990815, -5.8188143e-05, -2.9736952e-06, 0.0010021529, 0.00048666264, -6.131788e-05, -2.1386436e-06, 0.0012366746, 0.00045106385, -6.3900196e-05, -1.326115e-06, 0.0014528794, 0.00041345222, -6.5939574e-05, -5.401463e-07, 0.0016498462, 0.00037416894, -6.744375e-05, 2.155066e-07, 0.0018268245, 0.00033355382, -6.842356e-05, 9.3738475e-07, 0.0019832323, 0.00029194297, -6.889279e-05, 1.6223406e-06, 0.0021186548, 0.00024966677, -6.886801e-05, 2.2675495e-06, 0.0022328403, 0.00020704798, -6.836832e-05, 2.870518e-06, 0.0023256964, 0.00016439987, -6.741521e-05, 3.4290915e-06, 0.0023972844, 0.00012202443, -6.603233e-05, 3.941457e-06, 0.0024478133, 8.021083e-05, -6.4245236e-05, 4.4061467e-06, 0.0024776335, 3.923397e-05, -6.208121e-05, 4.822034e-06, 0.002487229, -6.469001e-07, -5.9569018e-05, 5.188334e-06, 0.0024772089, -3.918929e-05, -5.6738638e-05, 5.504596e-06, 0.0024482994, -7.616852e-05, -5.3621086e-05, 5.7706984e-06, 0.0024013345, -0.0001113786, -5.0248134e-05, 5.9868366e-06, 0.0023372462, -0.00014463293, -4.6652112e-05, 6.153516e-06, 0.0022570551, -0.00017576489, -4.2865657e-05, 6.271535e-06, 0.0021618593, -0.00020462825, -3.8921502e-05, 6.3419734e-06, 0.0020528259, -0.00023109744, -3.4852266e-05, 6.366177e-06, 0.0019311786, -0.0002550677, -3.069023e-05, 6.345739e-06, 0.0017981889, -0.00027645496, -2.6467147e-05, 6.2824834e-06, 0.0016551651, -0.00029519593, -2.221406e-05, 6.178445e-06, 0.0015034418, -0.00031124748, -1.7961107e-05, 6.03585e-06, 0.0013443704, -0.00032458652, -1.3737362e-05, 5.857096e-06, 0.0011793087, -0.00033520933, -9.570685e-06, 5.644729e-06, 0.0010096121, -0.00034313093, -5.48757e-06, 5.4014263e-06, 0.0008366235, -0.00034838438, -1.5130255e-06, 5.12997e-06, 0.0006616651, -0.00035101993, 2.3295459e-06, 4.8332295e-06, 0.00048602998, -0.00035110404, 6.0184434e-06, 4.514138e-06, 0.0003109739, -0.00034871852, 9.533757e-06, 4.1756716e-06, 0.00013770835, -0.00034395925, 1.2857436e-05, 3.8208295e-06, -3.260657e-05, -0.0003369353, 1.5973346e-05, 3.4526136e-06, -0.00019886826, -0.00032776754, 1.8867311e-05, 3.0740066e-06, -0.00036003732, -0.0003165875, 2.1527147e-05, 2.6879568e-06, -0.00051514246, -0.00030353622, 2.3942659e-05, 2.2973575e-06, -0.0006632851, -0.0002887628, 2.6105663e-05, 1.9050303e-06, -0.0008036428, -0.0002724232, 2.8009958e-05, 1.5137099e-06, -0.0009354727, -0.00025467912, 2.96513e-05, 1.1260281e-06, -0.001058114, -0.00023569637, 3.102738e-05, 7.445007e-07, -0.0011709894, -0.00021564393, 3.2137745e-05, 3.7151443e-07, -0.0012736067, -0.00019469253, 3.2983775e-05, 9.315632e-09, -0.0013655593, -0.0001730135, 3.3568576e-05, -3.399997e-07, -0.001446526, -0.00015077756, 3.3896933e-05, -6.7449474e-07, -0.0015162709, -0.00012815373, 3.3975193e-05, -9.923992e-07, -0.0015746417, -0.000105308165, 3.381119e-05, -1.2921158e-06, -0.0016215681, -8.240324e-05, 3.3414137e-05, -1.5722242e-06, -0.0016570602, -5.9596467e-05, 3.2794516e-05, -1.8314852e-06, -0.0016812052, -3.7039645e-05, 3.1963966e-05, -2.0688426e-06, -0.0016941648, -1.4878019e-05, 3.0935164e-05, -2.2834242e-06, -0.0016961712, 6.7504993e-06, 2.972171e-05, -2.4745411e-06, -0.001687524, 2.7716016e-05, 2.8338003e-05, -2.6416863e-06, -0.0016685852, 4.7897276e-05, 2.6799118e-05, -2.7845317e-06, -0.0016397756, 6.71822e-05, 2.5120677e-05, -2.9029245e-06, -0.001601569, 8.546832e-05, 2.3318733e-05, -2.9968828e-06, -0.0015544887, 0.0001026632, 2.1409647e-05, -3.0665883e-06, -0.001499101, 0.0001186847, 1.9409963e-05, -3.1123816e-06, -0.0014360112, 0.00013346122, 1.7336295e-05, -3.134753e-06, -0.0013658573, 0.00014693181, 1.5205208e-05, -3.1343338e-06, -0.0012893054, 0.00015904625, 1.30331155e-05, -3.11189e-06, -0.0012070436, 0.00016976509, 1.083617e-05, -3.0683095e-06, -0.0011197778, 0.00017905947, 8.630162e-06, -3.0045944e-06, -0.0010282248, 0.00018691104, 6.430425e-06, -2.9218488e-06, -0.00093310873, 0.00019331177, 4.2517527e-06, -2.8212694e-06, -0.00083515485, 0.00019826357, 2.1083124e-06, -2.7041333e-06, -0.00073508505, 0.00020177808, 1.3571504e-08, -2.571787e-06, -0.00063361326, 0.00020387616, -2.01977e-06, -2.425636e-06, -0.0005314405, 0.00020458754, -3.979839e-06, -2.2671322e-06, -0.000429251, 0.00020395032, -5.8556443e-06, -2.0977627e-06, -0.00032770785, 0.0002020104, -7.637118e-06, -1.9190397e-06, -0.00022744942, 0.00019882098, -9.3151575e-06, -1.7324882e-06, -0.00012908576, 0.00019444192, -1.088165e-05, -1.5396362e-06, -3.319544e-05, 0.00018893916, -1.2329501e-05, -1.3420041e-06, 5.9677324e-05, 0.00018238404, -1.3652642e-05, -1.1410947e-06, 0.0001490252, 0.00017485271, -1.4846045e-05, -9.3838355e-07, 0.00023438, 0.00016642542, -1.5905714e-05, -7.353101e-07, 0.00031531454, 0.00015718587, -1.6828686e-05, -5.3326926e-07, 0.0003914442, 0.0001472205, -1.7613016e-05, -3.3360325e-07, 0.0004624281, 0.00013661788, -1.825775e-05, -1.3759457e-07, 0.00052797014, 0.00012546804, -1.8762907e-05, 5.3540806e-08, 0.0005878194, 0.000113861744, -1.9129448e-05, 2.3865942e-07, 0.0006417703, 0.00010188999, -1.9359228e-05, 4.1669557e-07, 0.0006896629, 8.964328e-05, -1.945497e-05, 5.8666603e-07, 0.00073138205, 7.721108e-05, -1.9420208e-05, 7.476739e-07, 0.0007668571, 6.468125e-05, -1.925924e-05, 8.9891165e-07, 0.0007960607, 5.2139505e-05, -1.897707e-05, 1.0396641e-06, 0.0008190079, 3.9668917e-05, -1.8579363e-05, 1.1693096e-06, 0.0008357543, 2.7349433e-05, -1.8072376e-05, 1.2873218e-06, 0.0008463948, 1.5257455e-05, -1.7462895e-05, 1.3932693e-06, 0.00085106137, 3.465429e-06, -1.6758184e-05, 1.4868162e-06, 0.0008499212, -7.958501e-06, -1.5965908e-05, 1.567721e-06, 0.00084317446, -1.8950814e-05, -1.5094076e-05, 1.6358349e-06, 0.0008310518, -2.9452885e-05, -1.41509745e-05, 1.6911001e-06, 0.00081381196, -3.941123e-05, -1.3145104e-05, 1.733547e-06, 0.000791739, -4.8777674e-05, -1.2085113e-05, 1.7632915e-06, 0.0007651399, -5.7509533e-05, -1.0979736e-05, 1.780531e-06, 0.0007343413, -6.55697e-05, -9.837733e-06, 1.7855406e-06, 0.0006996873, -7.292672e-05, -8.66783e-06, 1.7786688e-06, 0.000661536, -7.955482e-05, -7.4786617e-06, 1.7603329e-06, 0.0006202573, -8.543389e-05, -6.278715e-06, 1.7310136e-06, 0.0005762294, -9.0549445e-05, -5.0762783e-06, 1.6912501e-06, 0.00052983663, -9.4892544e-05, -3.879393e-06, 1.6416344e-06, 0.00048146633, -9.8459655e-05, -2.6958062e-06, 1.5828055e-06, 0.0004315062, -0.00010125252, -1.5329299e-06, 1.515444e-06, 0.0003803419, -0.00010327796, -3.9780068e-07, 1.4402657e-06, 0.0003283544, -0.00010454768, 7.029545e-07, 1.3580162e-06, 0.00027591767, -0.00010507803, 1.7631493e-06, 1.2694644e-06, 0.0002233964, -0.000104889725, 2.7770657e-06, 1.1753968e-06, 0.00017114387, -0.00010400761, 3.7394766e-06, 1.0766122e-06, 0.000119499964, -0.00010246032, 4.6456653e-06, 9.739147e-07, 6.878938e-05, -0.00010027998, 5.4914403e-06, 8.681094e-07, 1.9319938e-05, -9.75019e-05, 6.273147e-06, 7.599964e-07, -2.8618902e-05, -9.4164185e-05, 6.987674e-06, 6.5036573e-07, -7.4757394e-05, -9.030746e-05, 7.632458e-06, 5.399922e-07, -0.00011884663, -8.597446e-05, 8.205479e-06, 4.2963086e-07, -0.00016065953, -8.1209706e-05, 8.705265e-06, 3.200127e-07, -0.00019999166, -7.6059136e-05, 9.130872e-06, 2.1184024e-07, -0.00023666184, -7.0569775e-05, 9.481884e-06, 1.05784046e-07, -0.00027051257, -6.4789354e-05, 9.758393e-06, 2.4790348e-09, -0.00030141036, -5.8766007e-05, 9.960987e-06, -9.747847e-08, -0.00032924578, -5.25479e-05, 1.0090722e-05, -1.9353354e-07, -0.00035393343, -4.6182937e-05, 1.0149107e-05, -2.8517502e-07, -0.0003754118, -3.971843e-05, 1.01380765e-05, -3.7193755e-07, -0.00039364272, -3.3200828e-05, 1.00599655e-05, -4.5340315e-07, -0.00040861103, -2.6675398e-05, 9.917479e-06, -5.292025e-07, -0.00042032383, -2.0185998e-05, 9.713662e-06, -5.990159e-07, -0.0004288098, -1.377481e-05, 9.45187e-06, -6.625737e-07, -0.00043411818, -7.482119e-06, 9.135737e-06, -7.196567e-07, -0.00043631782, -1.3461047e-06, 8.76914e-06, -7.7009565e-07, -0.0004354962, 4.5973434e-06, 8.356164e-06, -8.137711e-07, -0.00043175797, 1.0314791e-05, 7.901073e-06, -8.506124e-07, -0.00042522405, 1.5775404e-05, 7.408275e-06, -8.805967e-07, -0.00041602994, 2.0951069e-05, 6.8822806e-06, -9.0374743e-07, -0.0004043246, 2.5816487e-05, 6.32768e-06, -9.2013283e-07, -0.0003902688, 3.0349262e-05, 5.7491015e-06, -9.29864e-07, -0.00037403396, 3.452994e-05, 5.151186e-06, -9.330925e-07, -0.00035580026, 3.834207e-05, 4.53855e-06, -9.3000864e-07, -0.00033575553, 4.177218e-05, 3.915759e-06, -9.208383e-07, -0.00031409352, 4.4809796e-05, 3.287298e-06, -9.058407e-07, -0.00029101243, 4.7447415e-05, 2.6575433e-06, -8.853054e-07, -0.00026671359, 4.9680435e-05, 2.0307386e-06, -8.5954946e-07, -0.00024139979, 5.150712e-05, 1.4109692e-06, -8.2891455e-07, -0.00021527409, 5.29285e-05, 8.0214056e-07, -7.937636e-07, -0.00018853832, 5.394828e-05, 2.0795864e-07, -7.544779e-07, -0.00016139183, 5.457273e-05, -3.6808916e-07, -7.11454e-07, -0.00013403017, 5.4810556e-05, -9.2274973e-07, -6.6510034e-07, -0.000106644016, 5.4672768e-05, -1.4530185e-06, -6.158344e-07, -7.941797e-05, 5.4172517e-05, -1.9561512e-06, -5.6407947e-07, -5.2529547e-05, 5.3324966e-05, -2.4296744e-06, -5.102617e-07, -2.6148235e-05, 5.2147087e-05, -2.8713919e-06, -4.548072e-07, -4.3459195e-07, 5.065752e-05, -3.2793919e-06, -3.98139e-07, 2.4460505e-05, 4.8876384e-05, -3.6520496e-06, -3.4067463e-07, 4.839657e-05, 4.6825076e-05, -3.988029e-06, -2.8282327e-07, 7.124411e-05, 4.4526125e-05, -4.286282e-06, -2.2498338e-07, 9.288513e-05, 4.2002965e-05, -4.5460474e-06, -1.6754049e-07, 0.000113213544, 3.9279777e-05, -4.7668445e-06, -1.1086485e-07, 0.0001321355, 3.6381287e-05, -4.9484693e-06, -5.530961e-08, 0.0001495696, 3.333259e-05, -5.0909857e-06, -1.2089328e-09, 0.00016544708, 3.015898e-05, -5.1947163e-06, 5.1123564e-08, 0.0001797118, 2.6885746e-05, -5.2602327e-06, 1.0139626e-07, 0.00019232024, 2.3538034e-05, -5.2883424e-06, 1.4934076e-07, 0.00020324139, 2.0140666e-05, -5.280078e-06, 1.9471295e-07, 0.00021245652, 1.6717991e-05, -5.2366795e-06, 2.3729379e-07, 0.00021995897, 1.3293736e-05, -5.1595825e-06, 2.7688998e-07, 0.00022575368, 9.890868e-06, -5.0504004e-06, 3.133345e-07, 0.00022985693, 6.531465e-06, -4.9109085e-06, 3.464867e-07, 0.00023229577, 3.2365963e-06, -4.7430276e-06, 3.7623255e-07, 0.0002331075, 2.6217998e-08, -4.5488046e-06, 4.0248443e-07, 0.0002323391, -3.0809283e-06, -4.3303958e-06, 4.2518093e-07, 0.0002300466, -6.067399e-06, -4.0900504e-06, 4.4428631e-07, 0.00022629442, -8.9171235e-06, -3.830089e-06, 4.5979002e-07, 0.00022115464, -1.1615467e-05, -3.55289e-06, 4.7170587e-07, 0.0002147063, -1.4149281e-05, -3.2608677e-06, 4.800712e-07, 0.00020703467, -1.6506945e-05, -2.9564578e-06, 4.849459e-07, 0.00019823038, -1.8678391e-05, -2.6420998e-06, 4.8641107e-07, 0.00018838872, -2.0655125e-05, -2.3202201e-06, 4.845681e-07, 0.00017760885, -2.243023e-05, -1.9932165e-06, 4.79537e-07, 0.00016599298, -2.3998355e-05, -1.6634432e-06, 4.7145537e-07, 0.00015364564, -2.5355715e-05, -1.3331963e-06, 4.604766e-07, 0.0001406728, -2.6500053e-05, -1.0047005e-06, 4.4676844e-07, 0.00012718125, -2.7430606e-05, -6.800967e-07, 4.3051145e-07, 0.00011327776, -2.814807e-05, -3.6142993e-07, 4.1189733e-07, 9.9068406e-05, -2.8654538e-05, -5.063932e-08, 3.9112732e-07, 8.465788e-05, -2.8953451e-05, 2.504517e-07, 3.6841044e-07, 7.014883e-05, -2.9049519e-05, 5.4014373e-07, 3.43962e-07, 5.5641256e-05, -2.894866e-05, 8.168688e-07, 3.1800187e-07, 4.1231902e-05, -2.8657914e-05, 1.0791964e-06, 2.9075287e-07, 2.701373e-05, -2.8185364e-05, 1.3258388e-06, 2.6243913e-07, 1.3075422e-05, -2.7540045e-05, 1.5556549e-06, 2.3328468e-07, -4.990741e-07, -2.6731852e-05, 1.767653e-06, 2.0351189e-07, -1.3630962e-05, -2.577145e-05, 1.960993e-06, 1.7333998e-07, -2.6246944e-05, -2.4670173e-05, 2.134986e-06, 1.4298375e-07, -3.8279537e-05, -2.3439934e-05, 2.2890958e-06, 1.12652266e-07, -4.9667346e-05, -2.209312e-05, 2.422936e-06, 8.254759e-08, -6.035525e-05, -2.064249e-05, 2.536268e-06, 5.2863736e-08, -7.0294605e-05, -1.9101093e-05, 2.6289983e-06, 2.3785605e-08, -7.944332e-05, -1.7482154e-05, 2.701174e-06, -4.5119646e-09, -8.7765955e-05, -1.579899e-05, 2.7529782e-06, -3.1865028e-08, -9.523373e-05, -1.4064918e-05, 2.784724e-06, -5.812128e-08, -0.0001018245, -1.22931615e-05, 2.7968485e-06, -8.3140684e-08, -0.0001075227, -1.0496768e-05, 2.789906e-06, -1.0679602e-07, -0.000112319205, -8.688526e-06, 2.7645597e-06, -1.2897331e-07, -0.00011621124, -6.8808913e-06, 2.7215747e-06, -1.4957217e-07, -0.00011920213, -5.0859103e-06, 2.6618093e-06, -1.6850602e-07, -0.00012130112, -3.3151562e-06, 2.5862055e-06, -1.8570219e-07, -0.0001225231, -1.579664e-06, 2.4957812e-06, -2.0110203e-07, -0.00012288833, 1.10123274e-07, 2.3916202e-06, -2.1466073e-07, -0.00012242218, 1.7444061e-06, 2.274863e-06, -2.2634732e-07, -0.000121154655, 3.3140732e-06, 2.1466967e-06, -2.361443e-07, -0.000119120225, 4.8107395e-06, 2.008347e-06, -2.4404736e-07, -0.00011635732, 6.2267804e-06, 1.8610679e-06, -2.5006503e-07, -0.000112908, 7.555355e-06, 1.7061315e-06, -2.542181e-07, -0.00010881753, 8.790428e-06, 1.5448207e-06, -2.565392e-07, -0.00010413401, 9.926786e-06, 1.3784193e-06, -2.5707212e-07, -9.890792e-05, 1.0960043e-05, 1.2082031e-06, -2.558712e-07, -9.319174e-05, 1.1886642e-05, 1.0354325e-06, -2.530006e-07, -8.703951e-05, 1.2703855e-05, 8.6134395e-07, -2.4853352e-07, -8.050644e-05, 1.3409771e-05, 6.871426e-07, -2.4255152e-07, -7.364849e-05, 1.4003287e-05, 5.1399525e-07, -2.3514356e-07, -6.6521956e-05, 1.4484084e-05, 3.430241e-07, -2.2640532e-07, -5.9183138e-05, 1.4852606e-05, 1.7530024e-07, -2.1643822e-07, -5.1687897e-05, 1.5110034e-05, 1.1838454e-08, -2.0534864e-07, -4.409134e-05, 1.5258252e-05, -1.4640786e-07, -1.9324698e-07, -3.6447458e-05, 1.529981e-05, -2.9855102e-07, -1.8024683e-07, -2.8808818e-05, 1.5237888e-05, -4.4377282e-07, -1.6646412e-07, -2.1226233e-05, 1.5076257e-05, -5.8132787e-07, -1.5201623e-07};
	localparam real hb[0:1199] = {0.027848251, 7.863854e-05, -0.000102238904, -5.581651e-07, 0.027769677, 0.00023546736, -0.000101059166, -1.6659997e-06, 0.027612986, 0.000390961, -9.87138e-05, -2.7490748e-06, 0.027379066, 0.0005442468, -9.5228235e-05, -3.7924478e-06, 0.027069231, 0.0006944717, -9.0638314e-05, -4.7825465e-06, 0.026685225, 0.00084080873, -8.498945e-05, -5.7071875e-06, 0.026229188, 0.0009824634, -7.833585e-05, -6.5555873e-06, 0.025703654, 0.001118679, -7.073963e-05, -7.3183596e-06, 0.02511152, 0.0012487425, -6.227e-05, -7.98751e-06, 0.024456035, 0.0013719881, -5.300233e-05, -8.556417e-06, 0.023740761, 0.0014878028, -4.301732e-05, -9.01981e-06, 0.022969553, 0.0015956288, -3.240009e-05, -9.373733e-06, 0.022146536, 0.0016949669, -2.1239324e-05, -9.615509e-06, 0.021276066, 0.0017853795, -9.626397e-06, -9.743692e-06, 0.0203627, 0.0018664917, 2.3454697e-06, -9.758017e-06, 0.019411169, 0.0019379936, 1.4582022e-05, -9.659341e-06, 0.018426342, 0.0019996406, 2.698878e-05, -9.449581e-06, 0.017413195, 0.0020512538, 3.9471804e-05, -9.131647e-06, 0.016376775, 0.0020927207, 5.193842e-05, -8.709373e-06, 0.01532217, 0.0021239934, 6.429791e-05, -8.187441e-06, 0.014254476, 0.0021450883, 7.646218e-05, -7.5713097e-06, 0.013178764, 0.0021560842, 8.834636e-05, -6.8671284e-06, 0.01210005, 0.0021571212, 9.9869336e-05, -6.0816633e-06, 0.011023269, 0.0021483973, 0.00011095432, -5.2222153e-06, 0.009953238, 0.0021301666, 0.000121529265, -4.296539e-06, 0.008894636, 0.0021027357, 0.00013152728, -3.3127621e-06, 0.007851977, 0.0020664614, 0.000140887, -2.2793056e-06, 0.006829583, 0.0020217458, 0.00014955288, -1.2048044e-06, 0.005831566, 0.0019690336, 0.00015747549, -9.803153e-08, 0.004861804, 0.0019088082, 0.0001646116, 1.0321777e-06, 0.0039239265, 0.001841587, 0.00017092444, 2.176997e-06, 0.0030212952, 0.0017679174, 0.00017638376, 3.3276792e-06, 0.0021569917, 0.0016883726, 0.00018096587, 4.4756216e-06, 0.0013338061, 0.0016035473, 0.00018465356, 5.6124286e-06, 0.0005542263, 0.001514053, 0.0001874362, 6.7299707e-06, -0.00017956895, 0.0014205141, 0.00018930952, 7.820437e-06, -0.00086571515, 0.0013235628, 0.00019027547, 8.876385e-06, -0.0015026652, 0.0012238359, 0.00019034215, 9.890792e-06, -0.0020891905, 0.0011219693, 0.00018952347, 1.0857087e-05, -0.0026243792, 0.001018595, 0.00018783894, 1.176919e-05, -0.0031076341, 0.00091433653, 0.00018531342, 1.26215455e-05, -0.0035386665, 0.0008098057, 0.00018197673, 1.3409146e-05, -0.00391749, 0.00070559845, 0.0001778634, 1.4127555e-05, -0.0042444114, 0.0006022919, 0.00017301223, 1.477292e-05, -0.0045200214, 0.00050044095, 0.00016746596, 1.5341988e-05, -0.0047451803, 0.00040057558, 0.00016127084, 1.5832109e-05, -0.0049210084, 0.0003031979, 0.00015447625, 1.6241243e-05, -0.0050488687, 0.00020878005, 0.00014713424, 1.6567954e-05, -0.0051303525, 0.00011776187, 0.00013929917, 1.6811402e-05, -0.0051672626, 3.0549036e-05, 0.0001310272, 1.6971335e-05, -0.0051615955, -5.2488434e-05, 0.00012237595, 1.7048078e-05, -0.0051155235, -0.00013101756, 0.000113403985, 1.7042508e-05, -0.005031377, -0.00020474338, 0.00010417048, 1.6956043e-05, -0.0049116225, -0.00027340974, 9.473475e-05, 1.6790598e-05, -0.0047588455, -0.00033679965, 8.515589e-05, 1.6548585e-05, -0.0045757308, -0.00039473572, 7.549234e-05, 1.6232862e-05, -0.0043650414, -0.00044707974, 6.580157e-05, 1.5846703e-05, -0.0041295993, -0.0004937327, 5.6139706e-05, 1.539378e-05, -0.0038722672, -0.000534634, 4.656119e-05, 1.4878104e-05, -0.0035959282, -0.0005697608, 3.711847e-05, 1.4304009e-05, -0.003303467, -0.00059912674, 2.7861719e-05, 1.3676101e-05, -0.002997754, -0.00062278105, 1.8838567e-05, 1.2999224e-05, -0.002681625, -0.0006408069, 1.0093863e-05, 1.2278419e-05, -0.002357867, -0.0006533199, 1.6694551e-06, 1.1518884e-05, -0.0020292008, -0.00066046615, -6.395991e-06, 1.072594e-05, -0.0016982675, -0.0006624206, -1.4067155e-05, 9.904985e-06, -0.0013676136, -0.0006593847, -2.1312191e-05, 9.0614585e-06, -0.0010396786, -0.0006515847, -2.8102844e-05, 8.200804e-06, -0.0007167833, -0.00063926884, -3.441452e-05, 7.3284336e-06, -0.00040111947, -0.0006227055, -4.0226332e-05, 6.4496917e-06, -9.4740004e-05, -0.00060218055, -4.5521145e-05, 5.5698206e-06, 0.00020044901, -0.0005779951, -5.028556e-05, 4.6939313e-06, 0.0004826953, -0.0005504629, -5.4509896e-05, 3.826971e-06, 0.0007504061, -0.00051990815, -5.8188143e-05, 2.9736952e-06, 0.0010021529, -0.00048666264, -6.131788e-05, 2.1386436e-06, 0.0012366746, -0.00045106385, -6.3900196e-05, 1.326115e-06, 0.0014528794, -0.00041345222, -6.5939574e-05, 5.401463e-07, 0.0016498462, -0.00037416894, -6.744375e-05, -2.155066e-07, 0.0018268245, -0.00033355382, -6.842356e-05, -9.3738475e-07, 0.0019832323, -0.00029194297, -6.889279e-05, -1.6223406e-06, 0.0021186548, -0.00024966677, -6.886801e-05, -2.2675495e-06, 0.0022328403, -0.00020704798, -6.836832e-05, -2.870518e-06, 0.0023256964, -0.00016439987, -6.741521e-05, -3.4290915e-06, 0.0023972844, -0.00012202443, -6.603233e-05, -3.941457e-06, 0.0024478133, -8.021083e-05, -6.4245236e-05, -4.4061467e-06, 0.0024776335, -3.923397e-05, -6.208121e-05, -4.822034e-06, 0.002487229, 6.469001e-07, -5.9569018e-05, -5.188334e-06, 0.0024772089, 3.918929e-05, -5.6738638e-05, -5.504596e-06, 0.0024482994, 7.616852e-05, -5.3621086e-05, -5.7706984e-06, 0.0024013345, 0.0001113786, -5.0248134e-05, -5.9868366e-06, 0.0023372462, 0.00014463293, -4.6652112e-05, -6.153516e-06, 0.0022570551, 0.00017576489, -4.2865657e-05, -6.271535e-06, 0.0021618593, 0.00020462825, -3.8921502e-05, -6.3419734e-06, 0.0020528259, 0.00023109744, -3.4852266e-05, -6.366177e-06, 0.0019311786, 0.0002550677, -3.069023e-05, -6.345739e-06, 0.0017981889, 0.00027645496, -2.6467147e-05, -6.2824834e-06, 0.0016551651, 0.00029519593, -2.221406e-05, -6.178445e-06, 0.0015034418, 0.00031124748, -1.7961107e-05, -6.03585e-06, 0.0013443704, 0.00032458652, -1.3737362e-05, -5.857096e-06, 0.0011793087, 0.00033520933, -9.570685e-06, -5.644729e-06, 0.0010096121, 0.00034313093, -5.48757e-06, -5.4014263e-06, 0.0008366235, 0.00034838438, -1.5130255e-06, -5.12997e-06, 0.0006616651, 0.00035101993, 2.3295459e-06, -4.8332295e-06, 0.00048602998, 0.00035110404, 6.0184434e-06, -4.514138e-06, 0.0003109739, 0.00034871852, 9.533757e-06, -4.1756716e-06, 0.00013770835, 0.00034395925, 1.2857436e-05, -3.8208295e-06, -3.260657e-05, 0.0003369353, 1.5973346e-05, -3.4526136e-06, -0.00019886826, 0.00032776754, 1.8867311e-05, -3.0740066e-06, -0.00036003732, 0.0003165875, 2.1527147e-05, -2.6879568e-06, -0.00051514246, 0.00030353622, 2.3942659e-05, -2.2973575e-06, -0.0006632851, 0.0002887628, 2.6105663e-05, -1.9050303e-06, -0.0008036428, 0.0002724232, 2.8009958e-05, -1.5137099e-06, -0.0009354727, 0.00025467912, 2.96513e-05, -1.1260281e-06, -0.001058114, 0.00023569637, 3.102738e-05, -7.445007e-07, -0.0011709894, 0.00021564393, 3.2137745e-05, -3.7151443e-07, -0.0012736067, 0.00019469253, 3.2983775e-05, -9.315632e-09, -0.0013655593, 0.0001730135, 3.3568576e-05, 3.399997e-07, -0.001446526, 0.00015077756, 3.3896933e-05, 6.7449474e-07, -0.0015162709, 0.00012815373, 3.3975193e-05, 9.923992e-07, -0.0015746417, 0.000105308165, 3.381119e-05, 1.2921158e-06, -0.0016215681, 8.240324e-05, 3.3414137e-05, 1.5722242e-06, -0.0016570602, 5.9596467e-05, 3.2794516e-05, 1.8314852e-06, -0.0016812052, 3.7039645e-05, 3.1963966e-05, 2.0688426e-06, -0.0016941648, 1.4878019e-05, 3.0935164e-05, 2.2834242e-06, -0.0016961712, -6.7504993e-06, 2.972171e-05, 2.4745411e-06, -0.001687524, -2.7716016e-05, 2.8338003e-05, 2.6416863e-06, -0.0016685852, -4.7897276e-05, 2.6799118e-05, 2.7845317e-06, -0.0016397756, -6.71822e-05, 2.5120677e-05, 2.9029245e-06, -0.001601569, -8.546832e-05, 2.3318733e-05, 2.9968828e-06, -0.0015544887, -0.0001026632, 2.1409647e-05, 3.0665883e-06, -0.001499101, -0.0001186847, 1.9409963e-05, 3.1123816e-06, -0.0014360112, -0.00013346122, 1.7336295e-05, 3.134753e-06, -0.0013658573, -0.00014693181, 1.5205208e-05, 3.1343338e-06, -0.0012893054, -0.00015904625, 1.30331155e-05, 3.11189e-06, -0.0012070436, -0.00016976509, 1.083617e-05, 3.0683095e-06, -0.0011197778, -0.00017905947, 8.630162e-06, 3.0045944e-06, -0.0010282248, -0.00018691104, 6.430425e-06, 2.9218488e-06, -0.00093310873, -0.00019331177, 4.2517527e-06, 2.8212694e-06, -0.00083515485, -0.00019826357, 2.1083124e-06, 2.7041333e-06, -0.00073508505, -0.00020177808, 1.3571504e-08, 2.571787e-06, -0.00063361326, -0.00020387616, -2.01977e-06, 2.425636e-06, -0.0005314405, -0.00020458754, -3.979839e-06, 2.2671322e-06, -0.000429251, -0.00020395032, -5.8556443e-06, 2.0977627e-06, -0.00032770785, -0.0002020104, -7.637118e-06, 1.9190397e-06, -0.00022744942, -0.00019882098, -9.3151575e-06, 1.7324882e-06, -0.00012908576, -0.00019444192, -1.088165e-05, 1.5396362e-06, -3.319544e-05, -0.00018893916, -1.2329501e-05, 1.3420041e-06, 5.9677324e-05, -0.00018238404, -1.3652642e-05, 1.1410947e-06, 0.0001490252, -0.00017485271, -1.4846045e-05, 9.3838355e-07, 0.00023438, -0.00016642542, -1.5905714e-05, 7.353101e-07, 0.00031531454, -0.00015718587, -1.6828686e-05, 5.3326926e-07, 0.0003914442, -0.0001472205, -1.7613016e-05, 3.3360325e-07, 0.0004624281, -0.00013661788, -1.825775e-05, 1.3759457e-07, 0.00052797014, -0.00012546804, -1.8762907e-05, -5.3540806e-08, 0.0005878194, -0.000113861744, -1.9129448e-05, -2.3865942e-07, 0.0006417703, -0.00010188999, -1.9359228e-05, -4.1669557e-07, 0.0006896629, -8.964328e-05, -1.945497e-05, -5.8666603e-07, 0.00073138205, -7.721108e-05, -1.9420208e-05, -7.476739e-07, 0.0007668571, -6.468125e-05, -1.925924e-05, -8.9891165e-07, 0.0007960607, -5.2139505e-05, -1.897707e-05, -1.0396641e-06, 0.0008190079, -3.9668917e-05, -1.8579363e-05, -1.1693096e-06, 0.0008357543, -2.7349433e-05, -1.8072376e-05, -1.2873218e-06, 0.0008463948, -1.5257455e-05, -1.7462895e-05, -1.3932693e-06, 0.00085106137, -3.465429e-06, -1.6758184e-05, -1.4868162e-06, 0.0008499212, 7.958501e-06, -1.5965908e-05, -1.567721e-06, 0.00084317446, 1.8950814e-05, -1.5094076e-05, -1.6358349e-06, 0.0008310518, 2.9452885e-05, -1.41509745e-05, -1.6911001e-06, 0.00081381196, 3.941123e-05, -1.3145104e-05, -1.733547e-06, 0.000791739, 4.8777674e-05, -1.2085113e-05, -1.7632915e-06, 0.0007651399, 5.7509533e-05, -1.0979736e-05, -1.780531e-06, 0.0007343413, 6.55697e-05, -9.837733e-06, -1.7855406e-06, 0.0006996873, 7.292672e-05, -8.66783e-06, -1.7786688e-06, 0.000661536, 7.955482e-05, -7.4786617e-06, -1.7603329e-06, 0.0006202573, 8.543389e-05, -6.278715e-06, -1.7310136e-06, 0.0005762294, 9.0549445e-05, -5.0762783e-06, -1.6912501e-06, 0.00052983663, 9.4892544e-05, -3.879393e-06, -1.6416344e-06, 0.00048146633, 9.8459655e-05, -2.6958062e-06, -1.5828055e-06, 0.0004315062, 0.00010125252, -1.5329299e-06, -1.515444e-06, 0.0003803419, 0.00010327796, -3.9780068e-07, -1.4402657e-06, 0.0003283544, 0.00010454768, 7.029545e-07, -1.3580162e-06, 0.00027591767, 0.00010507803, 1.7631493e-06, -1.2694644e-06, 0.0002233964, 0.000104889725, 2.7770657e-06, -1.1753968e-06, 0.00017114387, 0.00010400761, 3.7394766e-06, -1.0766122e-06, 0.000119499964, 0.00010246032, 4.6456653e-06, -9.739147e-07, 6.878938e-05, 0.00010027998, 5.4914403e-06, -8.681094e-07, 1.9319938e-05, 9.75019e-05, 6.273147e-06, -7.599964e-07, -2.8618902e-05, 9.4164185e-05, 6.987674e-06, -6.5036573e-07, -7.4757394e-05, 9.030746e-05, 7.632458e-06, -5.399922e-07, -0.00011884663, 8.597446e-05, 8.205479e-06, -4.2963086e-07, -0.00016065953, 8.1209706e-05, 8.705265e-06, -3.200127e-07, -0.00019999166, 7.6059136e-05, 9.130872e-06, -2.1184024e-07, -0.00023666184, 7.0569775e-05, 9.481884e-06, -1.05784046e-07, -0.00027051257, 6.4789354e-05, 9.758393e-06, -2.4790348e-09, -0.00030141036, 5.8766007e-05, 9.960987e-06, 9.747847e-08, -0.00032924578, 5.25479e-05, 1.0090722e-05, 1.9353354e-07, -0.00035393343, 4.6182937e-05, 1.0149107e-05, 2.8517502e-07, -0.0003754118, 3.971843e-05, 1.01380765e-05, 3.7193755e-07, -0.00039364272, 3.3200828e-05, 1.00599655e-05, 4.5340315e-07, -0.00040861103, 2.6675398e-05, 9.917479e-06, 5.292025e-07, -0.00042032383, 2.0185998e-05, 9.713662e-06, 5.990159e-07, -0.0004288098, 1.377481e-05, 9.45187e-06, 6.625737e-07, -0.00043411818, 7.482119e-06, 9.135737e-06, 7.196567e-07, -0.00043631782, 1.3461047e-06, 8.76914e-06, 7.7009565e-07, -0.0004354962, -4.5973434e-06, 8.356164e-06, 8.137711e-07, -0.00043175797, -1.0314791e-05, 7.901073e-06, 8.506124e-07, -0.00042522405, -1.5775404e-05, 7.408275e-06, 8.805967e-07, -0.00041602994, -2.0951069e-05, 6.8822806e-06, 9.0374743e-07, -0.0004043246, -2.5816487e-05, 6.32768e-06, 9.2013283e-07, -0.0003902688, -3.0349262e-05, 5.7491015e-06, 9.29864e-07, -0.00037403396, -3.452994e-05, 5.151186e-06, 9.330925e-07, -0.00035580026, -3.834207e-05, 4.53855e-06, 9.3000864e-07, -0.00033575553, -4.177218e-05, 3.915759e-06, 9.208383e-07, -0.00031409352, -4.4809796e-05, 3.287298e-06, 9.058407e-07, -0.00029101243, -4.7447415e-05, 2.6575433e-06, 8.853054e-07, -0.00026671359, -4.9680435e-05, 2.0307386e-06, 8.5954946e-07, -0.00024139979, -5.150712e-05, 1.4109692e-06, 8.2891455e-07, -0.00021527409, -5.29285e-05, 8.0214056e-07, 7.937636e-07, -0.00018853832, -5.394828e-05, 2.0795864e-07, 7.544779e-07, -0.00016139183, -5.457273e-05, -3.6808916e-07, 7.11454e-07, -0.00013403017, -5.4810556e-05, -9.2274973e-07, 6.6510034e-07, -0.000106644016, -5.4672768e-05, -1.4530185e-06, 6.158344e-07, -7.941797e-05, -5.4172517e-05, -1.9561512e-06, 5.6407947e-07, -5.2529547e-05, -5.3324966e-05, -2.4296744e-06, 5.102617e-07, -2.6148235e-05, -5.2147087e-05, -2.8713919e-06, 4.548072e-07, -4.3459195e-07, -5.065752e-05, -3.2793919e-06, 3.98139e-07, 2.4460505e-05, -4.8876384e-05, -3.6520496e-06, 3.4067463e-07, 4.839657e-05, -4.6825076e-05, -3.988029e-06, 2.8282327e-07, 7.124411e-05, -4.4526125e-05, -4.286282e-06, 2.2498338e-07, 9.288513e-05, -4.2002965e-05, -4.5460474e-06, 1.6754049e-07, 0.000113213544, -3.9279777e-05, -4.7668445e-06, 1.1086485e-07, 0.0001321355, -3.6381287e-05, -4.9484693e-06, 5.530961e-08, 0.0001495696, -3.333259e-05, -5.0909857e-06, 1.2089328e-09, 0.00016544708, -3.015898e-05, -5.1947163e-06, -5.1123564e-08, 0.0001797118, -2.6885746e-05, -5.2602327e-06, -1.0139626e-07, 0.00019232024, -2.3538034e-05, -5.2883424e-06, -1.4934076e-07, 0.00020324139, -2.0140666e-05, -5.280078e-06, -1.9471295e-07, 0.00021245652, -1.6717991e-05, -5.2366795e-06, -2.3729379e-07, 0.00021995897, -1.3293736e-05, -5.1595825e-06, -2.7688998e-07, 0.00022575368, -9.890868e-06, -5.0504004e-06, -3.133345e-07, 0.00022985693, -6.531465e-06, -4.9109085e-06, -3.464867e-07, 0.00023229577, -3.2365963e-06, -4.7430276e-06, -3.7623255e-07, 0.0002331075, -2.6217998e-08, -4.5488046e-06, -4.0248443e-07, 0.0002323391, 3.0809283e-06, -4.3303958e-06, -4.2518093e-07, 0.0002300466, 6.067399e-06, -4.0900504e-06, -4.4428631e-07, 0.00022629442, 8.9171235e-06, -3.830089e-06, -4.5979002e-07, 0.00022115464, 1.1615467e-05, -3.55289e-06, -4.7170587e-07, 0.0002147063, 1.4149281e-05, -3.2608677e-06, -4.800712e-07, 0.00020703467, 1.6506945e-05, -2.9564578e-06, -4.849459e-07, 0.00019823038, 1.8678391e-05, -2.6420998e-06, -4.8641107e-07, 0.00018838872, 2.0655125e-05, -2.3202201e-06, -4.845681e-07, 0.00017760885, 2.243023e-05, -1.9932165e-06, -4.79537e-07, 0.00016599298, 2.3998355e-05, -1.6634432e-06, -4.7145537e-07, 0.00015364564, 2.5355715e-05, -1.3331963e-06, -4.604766e-07, 0.0001406728, 2.6500053e-05, -1.0047005e-06, -4.4676844e-07, 0.00012718125, 2.7430606e-05, -6.800967e-07, -4.3051145e-07, 0.00011327776, 2.814807e-05, -3.6142993e-07, -4.1189733e-07, 9.9068406e-05, 2.8654538e-05, -5.063932e-08, -3.9112732e-07, 8.465788e-05, 2.8953451e-05, 2.504517e-07, -3.6841044e-07, 7.014883e-05, 2.9049519e-05, 5.4014373e-07, -3.43962e-07, 5.5641256e-05, 2.894866e-05, 8.168688e-07, -3.1800187e-07, 4.1231902e-05, 2.8657914e-05, 1.0791964e-06, -2.9075287e-07, 2.701373e-05, 2.8185364e-05, 1.3258388e-06, -2.6243913e-07, 1.3075422e-05, 2.7540045e-05, 1.5556549e-06, -2.3328468e-07, -4.990741e-07, 2.6731852e-05, 1.767653e-06, -2.0351189e-07, -1.3630962e-05, 2.577145e-05, 1.960993e-06, -1.7333998e-07, -2.6246944e-05, 2.4670173e-05, 2.134986e-06, -1.4298375e-07, -3.8279537e-05, 2.3439934e-05, 2.2890958e-06, -1.12652266e-07, -4.9667346e-05, 2.209312e-05, 2.422936e-06, -8.254759e-08, -6.035525e-05, 2.064249e-05, 2.536268e-06, -5.2863736e-08, -7.0294605e-05, 1.9101093e-05, 2.6289983e-06, -2.3785605e-08, -7.944332e-05, 1.7482154e-05, 2.701174e-06, 4.5119646e-09, -8.7765955e-05, 1.579899e-05, 2.7529782e-06, 3.1865028e-08, -9.523373e-05, 1.4064918e-05, 2.784724e-06, 5.812128e-08, -0.0001018245, 1.22931615e-05, 2.7968485e-06, 8.3140684e-08, -0.0001075227, 1.0496768e-05, 2.789906e-06, 1.0679602e-07, -0.000112319205, 8.688526e-06, 2.7645597e-06, 1.2897331e-07, -0.00011621124, 6.8808913e-06, 2.7215747e-06, 1.4957217e-07, -0.00011920213, 5.0859103e-06, 2.6618093e-06, 1.6850602e-07, -0.00012130112, 3.3151562e-06, 2.5862055e-06, 1.8570219e-07, -0.0001225231, 1.579664e-06, 2.4957812e-06, 2.0110203e-07, -0.00012288833, -1.10123274e-07, 2.3916202e-06, 2.1466073e-07, -0.00012242218, -1.7444061e-06, 2.274863e-06, 2.2634732e-07, -0.000121154655, -3.3140732e-06, 2.1466967e-06, 2.361443e-07, -0.000119120225, -4.8107395e-06, 2.008347e-06, 2.4404736e-07, -0.00011635732, -6.2267804e-06, 1.8610679e-06, 2.5006503e-07, -0.000112908, -7.555355e-06, 1.7061315e-06, 2.542181e-07, -0.00010881753, -8.790428e-06, 1.5448207e-06, 2.565392e-07, -0.00010413401, -9.926786e-06, 1.3784193e-06, 2.5707212e-07, -9.890792e-05, -1.0960043e-05, 1.2082031e-06, 2.558712e-07, -9.319174e-05, -1.1886642e-05, 1.0354325e-06, 2.530006e-07, -8.703951e-05, -1.2703855e-05, 8.6134395e-07, 2.4853352e-07, -8.050644e-05, -1.3409771e-05, 6.871426e-07, 2.4255152e-07, -7.364849e-05, -1.4003287e-05, 5.1399525e-07, 2.3514356e-07, -6.6521956e-05, -1.4484084e-05, 3.430241e-07, 2.2640532e-07, -5.9183138e-05, -1.4852606e-05, 1.7530024e-07, 2.1643822e-07, -5.1687897e-05, -1.5110034e-05, 1.1838454e-08, 2.0534864e-07, -4.409134e-05, -1.5258252e-05, -1.4640786e-07, 1.9324698e-07, -3.6447458e-05, -1.529981e-05, -2.9855102e-07, 1.8024683e-07, -2.8808818e-05, -1.5237888e-05, -4.4377282e-07, 1.6646412e-07, -2.1226233e-05, -1.5076257e-05, -5.8132787e-07, 1.5201623e-07};
endpackage
`endif
