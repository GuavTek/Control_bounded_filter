`include "ComplexType.sv"

module RecursionModule #(
) (
    input complex in,
    output complex out
);
    
endmodule