`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam N = 4;
	localparam COEFF_BIAS = 48;
	localparam logic signed[63:0] Lfr[0:3] = {'d277489893271481, 'd277489893271481, 'd275315491622285, 'd275315491622285};
	localparam logic signed[63:0] Lfi[0:3] = {'d30020001337947, - 'd30020001337947, 'd11558098293529, - 'd11558098293529};
	localparam logic signed[63:0] Lbr[0:3] = {'d277489893271481, 'd277489893271481, 'd275315491622285, 'd275315491622285};
	localparam logic signed[63:0] Lbi[0:3] = {'d30020001337947, - 'd30020001337947, 'd11558098293529, - 'd11558098293529};
	localparam logic signed[63:0] Wfr[0:3] = {'d24193209882, 'd24193209882, - 'd7887428590, - 'd7887428590};
	localparam logic signed[63:0] Wfi[0:3] = {'d29297075841, - 'd29297075841, - 'd33126712469, 'd33126712469};
	localparam logic signed[63:0] Wbr[0:3] = {- 'd24193209882, - 'd24193209882, 'd7887428590, 'd7887428590};
	localparam logic signed[63:0] Wbi[0:3] = {- 'd29297075841, 'd29297075841, 'd33126712469, - 'd33126712469};
	localparam logic signed[63:0] Ffr[0:3][0:79] = '{
		'{'d2678910912348682, 'd1633669149297615, - 'd134405106412023, - 'd14489081406757, 'd3471761733289509, 'd1534935316807140, - 'd154547576200402, - 'd12167341321049, 'd4211153497515380, 'd1420087166233641, - 'd172563932222687, - 'd9743629047954, 'd4889422534499934, 'd1290723849399400, - 'd188281223922595, - 'd7247706595933, 'd5499740975037776, 'd1148585763351890, - 'd201556008143343, - 'd4709673588602, 'd6036181793402482, 'd995532040410431, - 'd212275515540637, - 'd2159613203878, 'd6493772333226378, 'd833517040657504, - 'd220358442413966, 'd372755769329, 'd6868535890318197, 'd664566135678268, - 'd225755365061278, 'd2858416831816, 'd7157521071022570, 'd490751075721102, - 'd228448778179966, 'd5269379888993, 'd7358818790936519, 'd314165232382821, - 'd228452763163329, 'd7578988059119, 'd7471566924126414, 'd136899005473061, - 'd225812296327788, 'd9762203913194, 'd7495942755766966, - 'd38984324020268, - 'd220602211106000, 'd11795872177577, 'd7433143529741519, - 'd211472022825834, - 'd212925832011491, 'd13658956252499, 'd7285355515665612, - 'd378624356972050, - 'd202913301681643, 'd15332746247078, 'd7055712145579892, - 'd538595822537850, - 'd190719625501872, 'd16801036599608, 'd6748241887867779, - 'd689654930258371, - 'd176522461172683, 'd18050271736293, 'd6367806633571694, - 'd830202339184127, - 'd160519683075600, 'd19069658617453, 'd5920031467125635, - 'd958787157130758, - 'd142926753400873, 'd19851245422781, 'd5411226778650929, - 'd1074121249927379, - 'd123973933701595, 'd20389966031699, 'd4848303747586724, - 'd1175091427164946, - 'd103903371822373, 'd20683650356549},
		'{'d2678910912348222, 'd1633669149297648, - 'd134405106412032, - 'd14489081406755, 'd3471761733289070, 'd1534935316807172, - 'd154547576200411, - 'd12167341321048, 'd4211153497514966, 'd1420087166233671, - 'd172563932222695, - 'd9743629047952, 'd4889422534499551, 'd1290723849399429, - 'd188281223922603, - 'd7247706595932, 'd5499740975037427, 'd1148585763351916, - 'd201556008143349, - 'd4709673588600, 'd6036181793402171, 'd995532040410455, - 'd212275515540643, - 'd2159613203877, 'd6493772333226108, 'd833517040657526, - 'd220358442413972, 'd372755769330, 'd6868535890317968, 'd664566135678286, - 'd225755365061283, 'd2858416831817, 'd7157521071022387, 'd490751075721118, - 'd228448778179969, 'd5269379888994, 'd7358818790936382, 'd314165232382833, - 'd228452763163332, 'd7578988059119, 'd7471566924126326, 'd136899005473070, - 'd225812296327790, 'd9762203913194, 'd7495942755766923, - 'd38984324020262, - 'd220602211106001, 'd11795872177577, 'd7433143529741523, - 'd211472022825831, - 'd212925832011491, 'd13658956252499, 'd7285355515665663, - 'd378624356972050, - 'd202913301681642, 'd15332746247078, 'd7055712145579987, - 'd538595822537854, - 'd190719625501870, 'd16801036599608, 'd6748241887867917, - 'd689654930258378, - 'd176522461172680, 'd18050271736292, 'd6367806633571872, - 'd830202339184137, - 'd160519683075597, 'd19069658617452, 'd5920031467125852, - 'd958787157130771, - 'd142926753400869, 'd19851245422781, 'd5411226778651180, - 'd1074121249927394, - 'd123973933701590, 'd20389966031698, 'd4848303747587006, - 'd1175091427164964, - 'd103903371822367, 'd20683650356548},
		'{- 'd2621464726625032, - 'd1601298142322358, 'd114277463862052, - 'd54557765512014, - 'd3402192470904109, - 'd1521613693668172, 'd101035526953527, - 'd52555428834631, - 'd4143075592769200, - 'd1441949887694716, 'd88125723066021, - 'd50522608463608, - 'd4844167648167600, - 'd1362478337710847, 'd75562184921028, - 'd48464973598293, - 'd5505606112696863, - 'd1283363101544773, 'd63357707642890, - 'd46388011318305, - 'd6127608592847788, - 'd1204760640672868, 'd51523776702445, - 'd44297022280332, - 'd6710469021379336, - 'd1126819797494854, 'd40070597533593, - 'd42197116997554, - 'd7254553845722606, - 'd1049681790049648, 'd29007126689070, - 'd40093212685504, - 'd7760298217955961, - 'd973480223457764, 'd18341104403946, - 'd37990030657633, - 'd8228202194534652, - 'd898341117369665, 'd8079088437780, - 'd35892094253348, - 'd8658826953596720, - 'd824382948694780, - 'd1773510931025, - 'd33803727280864, - 'd9052791037303526, - 'd751716708882984, - 'd11212394882364, - 'd31729052956814, - 'd9410766626308762, - 'd680445975029133, - 'd20234339123843, - 'd29671993324251, - 'd9733475853085184, - 'd610666994071677, - 'd28837156170190, - 'd27636269130411, - 'd10021687160474126, - 'd542468779358319, - 'd37019656947170, - 'd25625400145358, - 'd10276211711460314, - 'd475933218855185, - 'd44781611831263, - 'd23642705902492, - 'd10497899855813746, - 'd411135194280852, - 'd52123711232903, - 'd21691306841762, - 'd10687637658882664, - 'd348142710452834, - 'd59047525827614, - 'd19774125836360, - 'd10846343497467206, - 'd287017034141629, - 'd65555466535792, - 'd17893890083631, - 'd10974964727353150, - 'd227812841736200, - 'd71650744348225, - 'd16053133340965},
		'{- 'd2621464726623828, - 'd1601298142322414, 'd114277463862073, - 'd54557765512018, - 'd3402192470902937, - 'd1521613693668227, 'd101035526953548, - 'd52555428834635, - 'd4143075592768060, - 'd1441949887694769, 'd88125723066041, - 'd50522608463611, - 'd4844167648166494, - 'd1362478337710898, 'd75562184921047, - 'd48464973598296, - 'd5505606112695792, - 'd1283363101544822, 'd63357707642909, - 'd46388011318308, - 'd6127608592846752, - 'd1204760640672916, 'd51523776702463, - 'd44297022280336, - 'd6710469021378337, - 'd1126819797494900, 'd40070597533610, - 'd42197116997558, - 'd7254553845721645, - 'd1049681790049693, 'd29007126689086, - 'd40093212685508, - 'd7760298217955038, - 'd973480223457806, 'd18341104403961, - 'd37990030657636, - 'd8228202194533767, - 'd898341117369706, 'd8079088437795, - 'd35892094253351, - 'd8658826953595873, - 'd824382948694820, - 'd1773510931011, - 'd33803727280867, - 'd9052791037302716, - 'd751716708883021, - 'd11212394882350, - 'd31729052956816, - 'd9410766626307994, - 'd680445975029168, - 'd20234339123830, - 'd29671993324253, - 'd9733475853084454, - 'd610666994071711, - 'd28837156170178, - 'd27636269130413, - 'd10021687160473434, - 'd542468779358351, - 'd37019656947158, - 'd25625400145361, - 'd10276211711459662, - 'd475933218855215, - 'd44781611831252, - 'd23642705902494, - 'd10497899855813134, - 'd411135194280880, - 'd52123711232892, - 'd21691306841764, - 'd10687637658882086, - 'd348142710452861, - 'd59047525827604, - 'd19774125836362, - 'd10846343497466668, - 'd287017034141654, - 'd65555466535783, - 'd17893890083633, - 'd10974964727352650, - 'd227812841736223, - 'd71650744348217, - 'd16053133340967}};
	localparam logic signed[63:0] Ffi[0:3][0:79] = '{
		'{- 'd7789584925020542, 'd708887221199158, 'd206702748225345, - 'd19845819841343, - 'd7393588604643268, 'd873085743790186, 'd189441643064671, - 'd21110141804839, - 'd6918639246994867, 'd1024429359565470, 'd170276674079435, - 'd22108944360993, - 'd6371556198568730, 'd1161381434685642, 'd149461551191332, - 'd22835111110926, - 'd5759879607888508, 'd1282597644249564, 'd127264837936302, - 'd23284800600437, - 'd5091771080218742, 'd1386938313763277, 'd103966594132111, - 'd23457435961284, - 'd4375908801885497, 'd1473478185138040, 'd79854941677750, - 'd23355656937657, - 'd3621378440744956, 'd1541513537288885, 'd55222594523002, - 'd22985235482842, - 'd2837561156357778, 'd1590566623196748, 'd30363393574268, - 'd22354956512906, - 'd2034020064558232, 'd1620387416998140, 'd5568886563156, - 'd21476465781011, - 'd1220386496487038, 'd1630952695911008, - 'd18875008286193, - 'd20364087183631, - 'd406247372102465, 'd1622462512239921, - 'd42691217575166, - 'd19034612125145, 'd398965026813756, 'd1595334139989243, - 'd65614571842042, - 'd17507063846684, 'd1186079648425665, 'd1550193608429831, - 'd87394675671855, - 'd15802439866300, 'd1946288454422587, 'd1487864961015521, - 'd107798558746626, - 'd13943435878179, 'd2671242297735851, 'd1409357402058381, - 'd126613080816752, - 'd11954154617209, 'd3353139883456778, 'd1315850515302490, - 'd143647066875003, - 'd9859803310541, 'd3984808899006887, 'd1208677757771555, - 'd158733152334642, - 'd7686383409257, 'd4559778505553668, 'd1089308448825112, - 'd171729321708043, - 'd5460376320793, 'd5072342496187033, 'd959328488094488, - 'd182520128106280, - 'd3208428846785},
		'{'d7789584925020678, - 'd708887221199165, - 'd206702748225342, 'd19845819841342, 'd7393588604643451, - 'd873085743790196, - 'd189441643064668, 'd21110141804838, 'd6918639246995094, - 'd1024429359565484, - 'd170276674079431, 'd22108944360992, 'd6371556198568998, - 'd1161381434685658, - 'd149461551191327, 'd22835111110925, 'd5759879607888814, - 'd1282597644249583, - 'd127264837936296, 'd23284800600436, 'd5091771080219080, - 'd1386938313763298, - 'd103966594132105, 'd23457435961283, 'd4375908801885863, - 'd1473478185138064, - 'd79854941677743, 'd23355656937656, 'd3621378440745346, - 'd1541513537288910, - 'd55222594522994, 'd22985235482840, 'd2837561156358186, - 'd1590566623196775, - 'd30363393574260, 'd22354956512905, 'd2034020064558654, - 'd1620387416998168, - 'd5568886563148, 'd21476465781009, 'd1220386496487468, - 'd1630952695911038, 'd18875008286202, 'd20364087183629, 'd406247372102900, - 'd1622462512239951, 'd42691217575174, 'd19034612125143, - 'd398965026813322, - 'd1595334139989273, 'd65614571842050, 'd17507063846682, - 'd1186079648425238, - 'd1550193608429861, 'd87394675671863, 'd15802439866299, - 'd1946288454422172, - 'd1487864961015550, 'd107798558746634, 'd13943435878177, - 'd2671242297735452, - 'd1409357402058410, 'd126613080816760, 'd11954154617207, - 'd3353139883456400, - 'd1315850515302518, 'd143647066875011, 'd9859803310540, - 'd3984808899006532, - 'd1208677757771581, 'd158733152334649, 'd7686383409256, - 'd4559778505553342, - 'd1089308448825137, 'd171729321708049, 'd5460376320792, - 'd5072342496186738, - 'd959328488094511, 'd182520128106285, 'd3208428846784},
		'{'d20410122023596984, - 'd1087203619517777, 'd261581401330405, - 'd19688353631198, 'd19855845437227768, - 'd1129165953014674, 'd260549776479662, - 'd21497800075813, 'd19281639300793944, - 'd1166937977762846, 'd258996978016206, - 'd23185429430581, 'd18689575854732616, - 'd1200612237457261, 'd256948048973282, - 'd24752655664962, 'd18081679793730520, - 'd1230286297560720, 'd254428064696757, - 'd26201094598827, 'd17459925861202104, - 'd1256062325165291, 'd251462077212791, - 'd27532552007075, 'd16826236651983674, - 'd1278046676369314, 'd248075061960339, - 'd28749011807856, 'd16182480619338714, - 'd1296349491750649, 'd244291866905447, - 'd29852624356494, 'd15530470282089826, - 'd1311084300475151, 'd240137164048391, - 'd30845694866052, 'd14871960627433400, - 'd1322367633538259, 'd235635403329143, - 'd31730671974348, 'd14208647704754270, - 'd1330318646597064, 'd230810768931151, - 'd32510136476076, 'd13542167405539158, - 'd1335058752810478, 'd225687137978284, - 'd33186790237559, 'd12874094424288384, - 'd1336711266066034, 'd220288041614798, - 'd33763445310536, 'd12205941395145922, - 'd1335401054933668, 'd214636628453457, - 'd34243013260277, 'd11539158198806890, - 'd1331254207649389, 'd208755630372409, - 'd34628494722203, 'd10875131434119388, - 'd1324397708395326, 'd202667330637182, - 'd34922969200132, 'd10215184048673250, - 'd1314959125107046, 'd196393534320064, - 'd35129585118164, 'd9560575122561506, - 'd1303066309004502, 'd189955540985356, - 'd35251550137213, 'd8912499799410572, - 'd1288847106009427, 'd183374119605357, - 'd35292121746123, 'd8272089358702066, - 'd1272429080179444, 'd176669485668604, - 'd35254598136332},
		'{- 'd20410122023597112, 'd1087203619517783, - 'd261581401330408, 'd19688353631199, - 'd19855845437227944, 'd1129165953014683, - 'd260549776479665, 'd21497800075814, - 'd19281639300794168, 'd1166937977762856, - 'd258996978016210, 'd23185429430582, - 'd18689575854732880, 'd1200612237457274, - 'd256948048973287, 'd24752655664963, - 'd18081679793730820, 'd1230286297560734, - 'd254428064696763, 'd26201094598828, - 'd17459925861202444, 'd1256062325165307, - 'd251462077212797, 'd27532552007076, - 'd16826236651984046, 'd1278046676369332, - 'd248075061960346, 'd28749011807857, - 'd16182480619339120, 'd1296349491750668, - 'd244291866905454, 'd29852624356495, - 'd15530470282090264, 'd1311084300475172, - 'd240137164048399, 'd30845694866053, - 'd14871960627433864, 'd1322367633538281, - 'd235635403329152, 'd31730671974350, - 'd14208647704754760, 'd1330318646597088, - 'd230810768931160, 'd32510136476078, - 'd13542167405539672, 'd1335058752810502, - 'd225687137978293, 'd33186790237561, - 'd12874094424288920, 'd1336711266066060, - 'd220288041614808, 'd33763445310538, - 'd12205941395146478, 'd1335401054933694, - 'd214636628453467, 'd34243013260279, - 'd11539158198807466, 'd1331254207649416, - 'd208755630372419, 'd34628494722205, - 'd10875131434119980, 'd1324397708395354, - 'd202667330637193, 'd34922969200134, - 'd10215184048673856, 'd1314959125107074, - 'd196393534320075, 'd35129585118166, - 'd9560575122562122, 'd1303066309004531, - 'd189955540985367, 'd35251550137215, - 'd8912499799411199, 'd1288847106009456, - 'd183374119605368, 'd35292121746125, - 'd8272089358702702, 'd1272429080179473, - 'd176669485668615, 'd35254598136334}};
	localparam logic signed[63:0] Fbr[0:3][0:79] = '{
		'{- 'd2678910912348682, 'd1633669149297615, 'd134405106412023, - 'd14489081406757, - 'd3471761733289509, 'd1534935316807140, 'd154547576200402, - 'd12167341321049, - 'd4211153497515380, 'd1420087166233641, 'd172563932222687, - 'd9743629047954, - 'd4889422534499934, 'd1290723849399400, 'd188281223922595, - 'd7247706595933, - 'd5499740975037776, 'd1148585763351890, 'd201556008143343, - 'd4709673588602, - 'd6036181793402482, 'd995532040410431, 'd212275515540637, - 'd2159613203878, - 'd6493772333226378, 'd833517040657504, 'd220358442413966, 'd372755769329, - 'd6868535890318197, 'd664566135678268, 'd225755365061278, 'd2858416831816, - 'd7157521071022570, 'd490751075721102, 'd228448778179966, 'd5269379888993, - 'd7358818790936519, 'd314165232382821, 'd228452763163329, 'd7578988059119, - 'd7471566924126414, 'd136899005473061, 'd225812296327788, 'd9762203913194, - 'd7495942755766966, - 'd38984324020268, 'd220602211106000, 'd11795872177577, - 'd7433143529741519, - 'd211472022825834, 'd212925832011491, 'd13658956252499, - 'd7285355515665612, - 'd378624356972050, 'd202913301681643, 'd15332746247078, - 'd7055712145579892, - 'd538595822537850, 'd190719625501872, 'd16801036599608, - 'd6748241887867779, - 'd689654930258371, 'd176522461172683, 'd18050271736293, - 'd6367806633571694, - 'd830202339184127, 'd160519683075600, 'd19069658617453, - 'd5920031467125635, - 'd958787157130758, 'd142926753400873, 'd19851245422781, - 'd5411226778650929, - 'd1074121249927379, 'd123973933701595, 'd20389966031699, - 'd4848303747586724, - 'd1175091427164946, 'd103903371822373, 'd20683650356549},
		'{- 'd2678910912348222, 'd1633669149297648, 'd134405106412032, - 'd14489081406755, - 'd3471761733289070, 'd1534935316807172, 'd154547576200411, - 'd12167341321048, - 'd4211153497514966, 'd1420087166233671, 'd172563932222695, - 'd9743629047952, - 'd4889422534499551, 'd1290723849399429, 'd188281223922603, - 'd7247706595932, - 'd5499740975037427, 'd1148585763351916, 'd201556008143349, - 'd4709673588600, - 'd6036181793402171, 'd995532040410455, 'd212275515540643, - 'd2159613203877, - 'd6493772333226108, 'd833517040657526, 'd220358442413972, 'd372755769330, - 'd6868535890317968, 'd664566135678286, 'd225755365061283, 'd2858416831817, - 'd7157521071022387, 'd490751075721118, 'd228448778179969, 'd5269379888994, - 'd7358818790936382, 'd314165232382833, 'd228452763163332, 'd7578988059119, - 'd7471566924126326, 'd136899005473070, 'd225812296327790, 'd9762203913194, - 'd7495942755766923, - 'd38984324020262, 'd220602211106001, 'd11795872177577, - 'd7433143529741523, - 'd211472022825831, 'd212925832011491, 'd13658956252499, - 'd7285355515665663, - 'd378624356972050, 'd202913301681642, 'd15332746247078, - 'd7055712145579987, - 'd538595822537854, 'd190719625501870, 'd16801036599608, - 'd6748241887867917, - 'd689654930258378, 'd176522461172680, 'd18050271736292, - 'd6367806633571872, - 'd830202339184137, 'd160519683075597, 'd19069658617452, - 'd5920031467125852, - 'd958787157130771, 'd142926753400869, 'd19851245422781, - 'd5411226778651180, - 'd1074121249927394, 'd123973933701590, 'd20389966031698, - 'd4848303747587006, - 'd1175091427164964, 'd103903371822367, 'd20683650356548},
		'{'d2621464726625032, - 'd1601298142322358, - 'd114277463862052, - 'd54557765512014, 'd3402192470904109, - 'd1521613693668172, - 'd101035526953527, - 'd52555428834631, 'd4143075592769200, - 'd1441949887694716, - 'd88125723066021, - 'd50522608463608, 'd4844167648167600, - 'd1362478337710847, - 'd75562184921028, - 'd48464973598293, 'd5505606112696863, - 'd1283363101544773, - 'd63357707642890, - 'd46388011318305, 'd6127608592847788, - 'd1204760640672868, - 'd51523776702445, - 'd44297022280332, 'd6710469021379336, - 'd1126819797494854, - 'd40070597533593, - 'd42197116997554, 'd7254553845722606, - 'd1049681790049648, - 'd29007126689070, - 'd40093212685504, 'd7760298217955961, - 'd973480223457764, - 'd18341104403946, - 'd37990030657633, 'd8228202194534652, - 'd898341117369665, - 'd8079088437780, - 'd35892094253348, 'd8658826953596720, - 'd824382948694780, 'd1773510931025, - 'd33803727280864, 'd9052791037303526, - 'd751716708882984, 'd11212394882364, - 'd31729052956814, 'd9410766626308762, - 'd680445975029133, 'd20234339123843, - 'd29671993324251, 'd9733475853085184, - 'd610666994071677, 'd28837156170190, - 'd27636269130411, 'd10021687160474126, - 'd542468779358319, 'd37019656947170, - 'd25625400145358, 'd10276211711460314, - 'd475933218855185, 'd44781611831263, - 'd23642705902492, 'd10497899855813746, - 'd411135194280852, 'd52123711232903, - 'd21691306841762, 'd10687637658882664, - 'd348142710452834, 'd59047525827614, - 'd19774125836360, 'd10846343497467206, - 'd287017034141629, 'd65555466535792, - 'd17893890083631, 'd10974964727353150, - 'd227812841736200, 'd71650744348225, - 'd16053133340965},
		'{'d2621464726623828, - 'd1601298142322414, - 'd114277463862073, - 'd54557765512018, 'd3402192470902937, - 'd1521613693668227, - 'd101035526953548, - 'd52555428834635, 'd4143075592768060, - 'd1441949887694769, - 'd88125723066041, - 'd50522608463611, 'd4844167648166494, - 'd1362478337710898, - 'd75562184921047, - 'd48464973598296, 'd5505606112695792, - 'd1283363101544822, - 'd63357707642909, - 'd46388011318308, 'd6127608592846752, - 'd1204760640672916, - 'd51523776702463, - 'd44297022280336, 'd6710469021378337, - 'd1126819797494900, - 'd40070597533610, - 'd42197116997558, 'd7254553845721645, - 'd1049681790049693, - 'd29007126689086, - 'd40093212685508, 'd7760298217955038, - 'd973480223457806, - 'd18341104403961, - 'd37990030657636, 'd8228202194533767, - 'd898341117369706, - 'd8079088437795, - 'd35892094253351, 'd8658826953595873, - 'd824382948694820, 'd1773510931011, - 'd33803727280867, 'd9052791037302716, - 'd751716708883021, 'd11212394882350, - 'd31729052956816, 'd9410766626307994, - 'd680445975029168, 'd20234339123830, - 'd29671993324253, 'd9733475853084454, - 'd610666994071711, 'd28837156170178, - 'd27636269130413, 'd10021687160473434, - 'd542468779358351, 'd37019656947158, - 'd25625400145361, 'd10276211711459662, - 'd475933218855215, 'd44781611831252, - 'd23642705902494, 'd10497899855813134, - 'd411135194280880, 'd52123711232892, - 'd21691306841764, 'd10687637658882086, - 'd348142710452861, 'd59047525827604, - 'd19774125836362, 'd10846343497466668, - 'd287017034141654, 'd65555466535783, - 'd17893890083633, 'd10974964727352650, - 'd227812841736223, 'd71650744348217, - 'd16053133340967}};
	localparam logic signed[63:0] Fbi[0:3][0:79] = '{
		'{'d7789584925020542, 'd708887221199158, - 'd206702748225345, - 'd19845819841343, 'd7393588604643268, 'd873085743790186, - 'd189441643064671, - 'd21110141804839, 'd6918639246994867, 'd1024429359565470, - 'd170276674079435, - 'd22108944360993, 'd6371556198568730, 'd1161381434685642, - 'd149461551191332, - 'd22835111110926, 'd5759879607888508, 'd1282597644249564, - 'd127264837936302, - 'd23284800600437, 'd5091771080218742, 'd1386938313763277, - 'd103966594132111, - 'd23457435961284, 'd4375908801885497, 'd1473478185138040, - 'd79854941677750, - 'd23355656937657, 'd3621378440744956, 'd1541513537288885, - 'd55222594523002, - 'd22985235482842, 'd2837561156357778, 'd1590566623196748, - 'd30363393574268, - 'd22354956512906, 'd2034020064558232, 'd1620387416998140, - 'd5568886563156, - 'd21476465781011, 'd1220386496487038, 'd1630952695911008, 'd18875008286193, - 'd20364087183631, 'd406247372102465, 'd1622462512239921, 'd42691217575166, - 'd19034612125145, - 'd398965026813756, 'd1595334139989243, 'd65614571842042, - 'd17507063846684, - 'd1186079648425665, 'd1550193608429831, 'd87394675671855, - 'd15802439866300, - 'd1946288454422587, 'd1487864961015521, 'd107798558746626, - 'd13943435878179, - 'd2671242297735851, 'd1409357402058381, 'd126613080816752, - 'd11954154617209, - 'd3353139883456778, 'd1315850515302490, 'd143647066875003, - 'd9859803310541, - 'd3984808899006887, 'd1208677757771555, 'd158733152334642, - 'd7686383409257, - 'd4559778505553668, 'd1089308448825112, 'd171729321708043, - 'd5460376320793, - 'd5072342496187033, 'd959328488094488, 'd182520128106280, - 'd3208428846785},
		'{- 'd7789584925020678, - 'd708887221199165, 'd206702748225342, 'd19845819841342, - 'd7393588604643451, - 'd873085743790196, 'd189441643064668, 'd21110141804838, - 'd6918639246995094, - 'd1024429359565484, 'd170276674079431, 'd22108944360992, - 'd6371556198568998, - 'd1161381434685658, 'd149461551191327, 'd22835111110925, - 'd5759879607888814, - 'd1282597644249583, 'd127264837936296, 'd23284800600436, - 'd5091771080219080, - 'd1386938313763298, 'd103966594132105, 'd23457435961283, - 'd4375908801885863, - 'd1473478185138064, 'd79854941677743, 'd23355656937656, - 'd3621378440745346, - 'd1541513537288910, 'd55222594522994, 'd22985235482840, - 'd2837561156358186, - 'd1590566623196775, 'd30363393574260, 'd22354956512905, - 'd2034020064558654, - 'd1620387416998168, 'd5568886563148, 'd21476465781009, - 'd1220386496487468, - 'd1630952695911038, - 'd18875008286202, 'd20364087183629, - 'd406247372102900, - 'd1622462512239951, - 'd42691217575174, 'd19034612125143, 'd398965026813322, - 'd1595334139989273, - 'd65614571842050, 'd17507063846682, 'd1186079648425238, - 'd1550193608429861, - 'd87394675671863, 'd15802439866299, 'd1946288454422172, - 'd1487864961015550, - 'd107798558746634, 'd13943435878177, 'd2671242297735452, - 'd1409357402058410, - 'd126613080816760, 'd11954154617207, 'd3353139883456400, - 'd1315850515302518, - 'd143647066875011, 'd9859803310540, 'd3984808899006532, - 'd1208677757771581, - 'd158733152334649, 'd7686383409256, 'd4559778505553342, - 'd1089308448825137, - 'd171729321708049, 'd5460376320792, 'd5072342496186738, - 'd959328488094511, - 'd182520128106285, 'd3208428846784},
		'{- 'd20410122023596984, - 'd1087203619517777, - 'd261581401330405, - 'd19688353631198, - 'd19855845437227768, - 'd1129165953014674, - 'd260549776479662, - 'd21497800075813, - 'd19281639300793944, - 'd1166937977762846, - 'd258996978016206, - 'd23185429430581, - 'd18689575854732616, - 'd1200612237457261, - 'd256948048973282, - 'd24752655664962, - 'd18081679793730520, - 'd1230286297560720, - 'd254428064696757, - 'd26201094598827, - 'd17459925861202104, - 'd1256062325165291, - 'd251462077212791, - 'd27532552007075, - 'd16826236651983674, - 'd1278046676369314, - 'd248075061960339, - 'd28749011807856, - 'd16182480619338714, - 'd1296349491750649, - 'd244291866905447, - 'd29852624356494, - 'd15530470282089826, - 'd1311084300475151, - 'd240137164048391, - 'd30845694866052, - 'd14871960627433400, - 'd1322367633538259, - 'd235635403329143, - 'd31730671974348, - 'd14208647704754270, - 'd1330318646597064, - 'd230810768931151, - 'd32510136476076, - 'd13542167405539158, - 'd1335058752810478, - 'd225687137978284, - 'd33186790237559, - 'd12874094424288384, - 'd1336711266066034, - 'd220288041614798, - 'd33763445310536, - 'd12205941395145922, - 'd1335401054933668, - 'd214636628453457, - 'd34243013260277, - 'd11539158198806890, - 'd1331254207649389, - 'd208755630372409, - 'd34628494722203, - 'd10875131434119388, - 'd1324397708395326, - 'd202667330637182, - 'd34922969200132, - 'd10215184048673250, - 'd1314959125107046, - 'd196393534320064, - 'd35129585118164, - 'd9560575122561506, - 'd1303066309004502, - 'd189955540985356, - 'd35251550137213, - 'd8912499799410572, - 'd1288847106009427, - 'd183374119605357, - 'd35292121746123, - 'd8272089358702066, - 'd1272429080179444, - 'd176669485668604, - 'd35254598136332},
		'{'d20410122023597112, 'd1087203619517783, 'd261581401330408, 'd19688353631199, 'd19855845437227944, 'd1129165953014683, 'd260549776479665, 'd21497800075814, 'd19281639300794168, 'd1166937977762856, 'd258996978016210, 'd23185429430582, 'd18689575854732880, 'd1200612237457274, 'd256948048973287, 'd24752655664963, 'd18081679793730820, 'd1230286297560734, 'd254428064696763, 'd26201094598828, 'd17459925861202444, 'd1256062325165307, 'd251462077212797, 'd27532552007076, 'd16826236651984046, 'd1278046676369332, 'd248075061960346, 'd28749011807857, 'd16182480619339120, 'd1296349491750668, 'd244291866905454, 'd29852624356495, 'd15530470282090264, 'd1311084300475172, 'd240137164048399, 'd30845694866053, 'd14871960627433864, 'd1322367633538281, 'd235635403329152, 'd31730671974350, 'd14208647704754760, 'd1330318646597088, 'd230810768931160, 'd32510136476078, 'd13542167405539672, 'd1335058752810502, 'd225687137978293, 'd33186790237561, 'd12874094424288920, 'd1336711266066060, 'd220288041614808, 'd33763445310538, 'd12205941395146478, 'd1335401054933694, 'd214636628453467, 'd34243013260279, 'd11539158198807466, 'd1331254207649416, 'd208755630372419, 'd34628494722205, 'd10875131434119980, 'd1324397708395354, 'd202667330637193, 'd34922969200134, 'd10215184048673856, 'd1314959125107074, 'd196393534320075, 'd35129585118166, 'd9560575122562122, 'd1303066309004531, 'd189955540985367, 'd35251550137215, 'd8912499799411199, 'd1288847106009456, 'd183374119605368, 'd35292121746125, 'd8272089358702702, 'd1272429080179473, 'd176669485668615, 'd35254598136334}};
	localparam logic signed[63:0] hf[0:1999] = {'d7033096503296, - 'd32897980416, - 'd10967230464, 'd63928604, 'd7000245665792, - 'd98394423296, - 'd10337267712, 'd188110032, 'd6934845456384, - 'd162997501952, - 'd9086782464, 'd301512896, 'd6837488844800, - 'd226124627968, - 'd7233756672, 'd397524544, 'd6709056110592, - 'd287210536960, - 'd4804252672, 'd470098240, 'd6550703833088, - 'd345713672192, - 'd1831931776, 'd513814560, 'd6363853881344, - 'd401122131968, 'd1642511488, 'd523933696, 'd6150172966912, - 'd452959338496, 'd5571985920, 'd496438560, 'd5911558488064, - 'd500788854784, 'd9903706112, 'd428068320, 'd5650113888256, - 'd544219168768, 'd14579948544, 'd316342016, 'd5368126111744, - 'd582907527168, 'd19538849792, 'd159572240, 'd5068042010624, - 'd616563212288, 'd24715249664, - 'd43130884, 'd4752438460416, - 'd644950327296, 'd30041542656, - 'd291865696, 'd4423997194240, - 'd667889827840, 'd35448557568, - 'd585954240, 'd4085474918400, - 'd685260537856, 'd40866439168, - 'd923966848, 'd3739673690112, - 'd697000263680, 'd46225510400, - 'd1303755136, 'd3389412343808, - 'd703105531904, 'd51457126400, - 'd1722493184, 'd3037497131008, - 'd703630671872, 'd56494514176, - 'd2176726784, 'd2686692360192, - 'd698686832640, 'd61273546752, - 'd2662427904, 'd2339693658112, - 'd688439820288, 'd65733513216, - 'd3175056896, 'd1999099920384, - 'd673107279872, 'd69817778176, - 'd3709628672, 'd1667389456384, - 'd652956008448, 'd73474457600, - 'd4260784384, 'd1346895216640, - 'd628297957376, 'd76656959488, - 'd4822863872, 'd1039784017920, - 'd599486234624, 'd79324479488, - 'd5389984768, 'd748036685824, - 'd566910648320, 'd81442447360, - 'd5956117504, 'd473431015424, - 'd530992660480, 'd82982838272, - 'd6515166720, 'd217527091200, - 'd492180406272, 'd83924451328, - 'd7061048320, - 'd18344486912, - 'd450943287296, 'd84253073408, - 'd7587765248, - 'd233092038656, - 'd407766368256, 'd83961561088, - 'd8089484800, - 'd425869180928, - 'd363144806400, 'd83049857024, - 'd8560607232, - 'd596078428160, - 'd317578280960, 'd81524924416, - 'd8995835904, - 'd743372095488, - 'd271565209600, 'd79400542208, - 'd9390236672, - 'd867650306048, - 'd225597456384, 'd76697108480, - 'd9739302912, - 'd969056190464, - 'd180154810368, 'd73441320960, - 'd10038998016, - 'd1047968874496, - 'd135700045824, 'd69665783808, - 'd10285808640, - 'd1104993583104, - 'd92673966080, 'd65408569344, - 'd10476781568, - 'd1140949254144, - 'd51490967552, 'd60712722432, - 'd10609551360, - 'd1156854972416, - 'd12534914048, 'd55625695232, - 'd10682369024, - 'd1153913061376, 'd23844581376, 'd50198769664, - 'd10694119424, - 'd1133491388416, 'd57335398400, 'd44486422528, - 'd10644324352, - 'd1097103966208, 'd87665672192, 'd38545653760, - 'd10533150720, - 'd1046390308864, 'd114606071808, 'd32435316736, - 'd10361399296, - 'd983093477376, 'd137971515392, 'd26215440384, - 'd10130492416, - 'd909037731840, 'd157622370304, 'd19946518528, - 'd9842454528, - 'd826105724928, 'd173465124864, 'd13688829952, - 'd9499883520, - 'd736215171072, 'd185452544000, 'd7501764608, - 'd9105917952, - 'd641296105472, 'd193583169536, 'd1443165440, - 'd8664196096, - 'd543267749888, 'd197900484608, - 'd4431298048, - 'd8178812416, - 'd444016885760, 'd198491455488, - 'd10068722688, - 'd7654265856, - 'd345376227328, 'd195484614656, - 'd15419525120, - 'd7095408640, - 'd249104269312, 'd189047783424, - 'd20437946368, - 'd6507388928, - 'd156866412544, 'd179385237504, - 'd25082505216, - 'd5895589888, - 'd70217392128, 'd166734675968, - 'd29316399104, - 'd5265568768, 'd9414508544, 'd151363747840, - 'd33107843072, - 'd4622995968, 'd80741564416, 'd133566259200, - 'd36430344192, - 'd3973589248, 'd142628683776, 'd113658347520, - 'd39262916608, - 'd3323052544, 'd194103558144, 'd91974221824, - 'd41590218752, - 'd2677014272, 'd234364616704, 'd68861943808, - 'd43402641408, - 'd2040966400, 'd262786842624, 'd44679032832, - 'd44696309760, - 'd1420208256, 'd278925475840, 'd19788113920, - 'd45473042432, - 'd819790720, 'd282517438464, - 'd5447470592, - 'd45740224512, - 'd244465792, 'd273480531968, - 'd30667960320, - 'd45510623232, 'd301360416, 'd251910750208, - 'd55521345536, - 'd44802162688, 'd813669824, 'd218077265920, - 'd79667380224, - 'd43637624832, 'd1288869760, 'd172415664128, - 'd102781378560, - 'd42044309504, 'd1723824640, 'd115519225856, - 'd124557795328, - 'd40053633024, 'd2115882240, 'd48128520192, - 'd144713433088, - 'd37700722688, 'd2462894336, - 'd28880474112, - 'd162990424064, - 'd35023921152, 'd2763230464, - 'd114509742080, - 'd179158859776, - 'd32064319488, 'd3015787008, - 'd207653748736, - 'd193018920960, - 'd28865234944, 'd3219988736, - 'd307115032576, - 'd204402835456, - 'd25471664128, 'd3375784960, - 'd411620442112, - 'd213176172544, - 'd21929756672, 'd3483641344, - 'd519838269440, - 'd219238973440, - 'd18286260224, 'd3544522240, - 'd630395568128, - 'd222526259200, - 'd14587981824, 'd3559872512, - 'd741895634944, - 'd223008227328, - 'd10881244160, 'd3531590144, - 'd852935704576, - 'd220690022400, - 'd7211374080, 'd3461996544, - 'd962124054528, - 'd215611097088, - 'd3622200320, 'd3353801728, - 'd1068097273856, - 'd207844130816, - 'd155578656, 'd3210066176, - 'd1169536057344, - 'd197493669888, 'd3149049344, 'd3034159104, - 'd1265181130752, - 'd184694308864, 'd6255063040, 'd2829713920, - 'd1353847668736, - 'd169608675328, 'd9129030656, 'd2600581376, - 'd1434438467584, - 'd152425005056, 'd11741032448, 'd2350781696, - 'd1505956593664, - 'd133354577920, 'd14064936960, 'd2084455552, - 'd1567515475968, - 'd112628752384, 'd16078633984, 'd1805813376, - 'd1618349129728, - 'd90496016384, 'd17764208640, 'd1519086592, - 'd1657819234304, - 'd67218747392, 'd19108071424, 'd1228478592, - 'd1685421162496, - 'd43069902848, 'd20101029888, 'd938116672, - 'd1700789092352, - 'd18329671680, 'd20738314240, 'd652006464, - 'd1703698104320, 'd6717959680, 'd21019545600, 'd373988160, - 'd1694065885184, 'd31788576768, 'd20948656128, 'd107695488, - 'd1671951417344, 'd56600698880, 'd20533766144, - 'd143481952, - 'd1637553012736, 'd80879017984, 'd19787003904, - 'd376432992, - 'd1591204642816, 'd104357543936, 'd18724286464, - 'd588355264, - 'd1533370171392, 'd126782562304, 'd17365071872, - 'd776781440, - 'd1464636669952, 'd147915423744, 'd15732052992, - 'd939601280, - 'd1385706160128, 'd167535099904, 'd13850836992, - 'd1075078784, - 'd1297386569728, 'd185440518144, 'd11749591040, - 'd1181864704, - 'd1200580722688, 'd201452535808, 'd9458661376, - 'd1259004928, - 'd1096275197952, 'd215415816192, 'd7010174464, - 'd1305943424, - 'd985527877632, 'd227200188416, 'd4437632000, - 'd1322520576, - 'd869455364096, 'd236701794304, 'd1775485824, - 'd1308967168, - 'd749219348480, 'd243843940352, - 'd941283776, - 'd1265894400, - 'd626012913664, 'd248577572864, - 'd3677590016, - 'd1194278144, - 'd501046935552, 'd250881425408, - 'd6398656512, - 'd1095440768, - 'd375535730688, 'd250761838592, - 'd9070423040, - 'd971028672, - 'd250683834368, 'd248252301312, - 'd11659934720, - 'd822986240, - 'd127672295424, 'd243412647936, - 'd14135713792, - 'd653526912, - 'd7645917696, 'd236328009728, - 'd16468104192, - 'd465101920, 'd108299083776, 'd227107389440, - 'd18629595136, - 'd260366176, 'd219126661120, 'd215882104832, - 'd20595109888, - 'd42143052, 'd323871637504, 'd202803920896, - 'd22342254592, 'd186612704, 'd421649350656, 'd188043018240, - 'd23851552768, 'd422852640, 'd511664455680, 'd171785748480, - 'd25106614272, 'd663472896, 'd593218240512, 'd154232242176, - 'd26094284800, 'd905352320, 'd665715081216, 'd135593918464, - 'd26804754432, 'd1145390336, 'd728667193344, 'd116090904576, - 'd27231608832, 'd1380543744, 'd781698727936, 'd95949373440, - 'd27371864064, 'd1607862400, 'd824547606528, 'd75398856704, - 'd27225939968, 'd1824522752, 'd857067028480, 'd54669598720, - 'd26797602816, 'd2027859968, 'd879224750080, 'd33989888000, - 'd26093875200, 'd2215397376, 'd891101773824, 'd13583513600, - 'd25124898816, 'd2384873216, 'd892889333760, - 'd6332733440, - 'd23903772672, 'd2534263552, 'd884884701184, - 'd25551407104, - 'd22446352384, 'd2661804288, 'd867486269440, - 'd43876618240, - 'd20771020800, 'd2766007296, 'd841186934784, - 'd61126078464, - 'd18898444288, 'd2845674240, 'd806566887424, - 'd77132947456, - 'd16851289088, 'd2899907328, 'd764285681664, - 'd91747483648, - 'd14653930496, 'd2928114688, 'd715073060864, - 'd104838455296, - 'd12332148736, 'd2930013696, 'd659719585792, - 'd116294311936, - 'd9912799232, 'd2905629696, 'd599066345472, - 'd126024146944, - 'd7423496704, 'd2855291904, 'd533994668032, - 'd133958361088, - 'd4892274176, 'd2779624704, 'd465415241728, - 'd140049088512, - 'd2347257600, 'd2679536640, 'd394257203200, - 'd144270393344, 'd183660272, 'd2556206336, 'd321457225728, - 'd146618138624, 'd2673139712, 'd2411064576, 'd247948623872, - 'd147109675008, 'd5094700032, 'd2245774336, 'd174650785792, - 'd145783259136, 'd7423012352, 'd2062207744, 'd102458908672, - 'd142697250816, 'd9634170880, 'd1862423296, 'd32234213376, - 'd137929080832, 'd11705949184, 'd1648637312, - 'd35205341184, - 'd131574038528, 'd13618027520, 'd1423197824, - 'd99093577728, - 'd123743797248, 'd15352196096, 'd1188554880, - 'd158723964928, - 'd114564939776, 'd16892532736, 'd947231424, - 'd213456617472, - 'd104177123328, 'd18225549312, 'd701792896, - 'd262724354048, - 'd92731334656, 'd19340306432, 'd454817568, - 'd306037915648, - 'd80387866624, 'd20228497408, 'd208866800, - 'd342990127104, - 'd67314339840, 'd20884506624, - 'd33544018, - 'd373259010048, - 'd53683642368, 'd21305427968, - 'd269973504, - 'd396609880064, - 'd39671808000, 'd21491048448, - 'd498081024, - 'd412896460800, - 'd25455941632, 'd21443817472, - 'd715651776, - 'd422060851200, - 'd11212149760, 'd21168769024, - 'd920620160, - 'd424132542464, 'd2886491648, 'd20673421312, - 'd1111091072, - 'd419226353664, 'd16671883264, 'd19967651840, - 'd1285358592, - 'd407539548160, 'd29982767104, 'd19063545856, - 'd1441922816, - 'd389347966976, 'd42666471424, 'd17975222272, - 'd1579503232, - 'd365001244672, 'd54580543488, 'd16718628864, - 'd1697049984, - 'd334917435392, 'd65594208256, 'd15311344640, - 'd1793752448, - 'd299576754176, 'd75589697536, 'd13772339200, - 'd1869043840, - 'd259514777600, 'd84463378432, 'd12121732096, - 'd1922604416, - 'd215315218432, 'd92126724096, 'd10380551168, - 'd1954360704, - 'd167602061312, 'd98507071488, 'd8570467840, - 'd1964482176, - 'd117031575552, 'd103548190720, 'd6713540096, - 'd1953375744, - 'd64283930624, 'd107210645504, 'd4831954432, - 'd1921676416, - 'd10054776832, 'd109471981568, 'd2947766016, - 'd1870237312, 'd44953247744, 'd110326685696, 'd1082651264, - 'd1800114816, 'd100038934528, 'd109785948160, - 'd742337920, - 'd1712554752, 'd154510770176, 'd107877253120, - 'd2507003392, - 'd1608973312, 'd207694921728, 'd104643788800, - 'd4192218624, - 'd1490939392, 'd258942943232, 'd100143644672, - 'd5780130304, - 'd1360152832, 'd307638960128, 'd94448910336, - 'd7254341120, - 'd1218423808, 'd353206403072, 'd87644585984, - 'd8600073216, - 'd1067649472, 'd395114184704, 'd79827378176, - 'd9804311552, - 'd909791232, 'd432882253824, 'd71104356352, - 'd10855919616, - 'd746850816, 'd466086363136, 'd61591547904, - 'd11745739776, - 'd580847104, 'd494362230784, 'd51412426752, - 'd12466658304, - 'd413792224, 'd517408784384, 'd40696356864, - 'd13013656576, - 'd247669072, 'd534990848000, 'd29576974336, - 'd13383830528, - 'd84408840, 'd546940780544, 'd18190557184, - 'd13576387584, 'd74130096, 'd553159360512, 'd6674405888, - 'd13592614912, 'd226182256, 'd553615949824, - 'd4834780672, - 'd13435834368, 'd370093632, 'd548347740160, - 'd16202491904, - 'd13111324672, 'd504338656, 'd537458442240, - 'd27297931264, - 'd12626223104, 'd627535488, 'd521115828224, - 'd37995479040, - 'd11989416960, 'd738459264, 'd499548880896, - 'd48176078848, - 'd11211404288, 'd836053504, 'd473044221952, - 'd57728499712, - 'd10304146432, 'd919438912, 'd441941950464, - 'd66550517760, - 'd9280902144, 'd987920768, 'd406630694912, - 'd74549952512, - 'd8156052992, 'd1040993088, 'd367542566912, - 'd81645584384, - 'd6944914944, 'd1078341504, 'd325147328512, - 'd87767891968, - 'd5663543808, 'd1099843200, 'd279946461184, - 'd92859727872, - 'd4328539136, 'd1105564672, 'd232466825216, - 'd96876699648, - 'd2956838144, 'd1095757824, 'd183254220800, - 'd99787579392, - 'd1565513600, 'd1070853440, 'd132866760704, - 'd101574352896, - 'd171574784, 'd1031453312, 'd81868210176, - 'd102232301568, 'd1208231424, 'd978319616, 'd30821447680, - 'd101769781248, 'd2557609472, 'd912363520, - 'd19718068224, - 'd100207943680, 'd3860898560, 'd834631680, - 'd69208547328, - 'd97580294144, 'd5103242240, 'd746291840, - 'd117127929856, - 'd93932068864, 'd6270749696, 'd648616768, - 'd162979545088, - 'd89319563264, 'd7350639104, 'd542967744, - 'd206297481216, - 'd83809280000, 'd8331369472, 'd430777056, - 'd246651437056, - 'd77476986880, 'd9202753536, 'd313529888, - 'd283651080192, - 'd70406725632, 'd9956050944, 'd192746128, - 'd316949954560, - 'd62689660928, 'd10584052736, 'd69961976, - 'd346248708096, - 'd54422949888, 'd11081128960, - 'd53288364, - 'd371297878016, - 'd45708509184, 'd11443279872, - 'd175490560, - 'd391899774976, - 'd36651757568, 'd11668144128, - 'd295167552, - 'd407910121472, - 'd27360344064, 'd11755006976, - 'd410896192, - 'd419238739968, - 'd17942872064, 'd11704777728, - 'd521323040, - 'd425849716736, - 'd8507630592, 'd11519951872, - 'd625179008, - 'd427760877568, 'd838650880, 'd11204558848, - 'd721292672, - 'd425042903040, 'd9992007680, 'd10764085248, - 'd808602688, - 'd417817427968, 'd18852395008, 'd10205391872, - 'd886167872, - 'd406254944256, 'd27324768256, 'd9536608256, - 'd953176704, - 'd390571982848, 'd35320111104, 'd8767017984, - 'd1008954368, - 'd371027836928, 'd42756349952, 'd7906931200, - 'd1052968640, - 'd347921055744, 'd49559191552, 'd6967550976, - 'd1084833536, - 'd321585086464, 'd55662837760, 'd5960825344, - 'd1104311424, - 'd292384145408, 'd61010624512, 'd4899297280, - 'd1111313664, - 'd260708253696, 'd65555509248, 'd3795950592, - 'd1105899136, - 'd226968616960, 'd69260451840, 'd2664050688, - 'd1088270976, - 'd191592300544, 'd72098676736, 'd1516986752, - 'd1058772032, - 'd155017199616, 'd74053804032, 'd368114528, - 'd1017878592, - 'd117686788096, 'd75119886336, - 'd769398208, - 'd966192896, - 'd80044908544, 'd75301273600, - 'd1882721152, - 'd904433792, - 'd42530721792, 'd74612400128, - 'd2959504384, - 'd833426688, - 'd5573702144, 'd73077473280, - 'd3988013824, - 'd754092160, 'd30411114496, 'd70729965568, - 'd4957257216, - 'd667433984, 'd65027657728, 'd67612160000, - 'd5857098752, - 'd574525888, 'd97903050752, 'd63774429184, - 'd6678363136, - 'd476498048, 'd128691486720, 'd59274575872, - 'd7412924928, - 'd374523168, 'd157077749760, 'd54177009664, - 'd8053787136, - 'd269802144, 'd182780313600, 'd48551907328, - 'd8595142656, - 'd163549664, 'd205553975296, 'd42474287104, - 'd9032420352, - 'd56980000, 'd225192067072, 'd36023083008, - 'd9362321408, 'd48707084, 'd241528176640, 'd29280149504, - 'd9582834688, 'd152339968, 'd254437326848, 'd22329272320, - 'd9693236224, 'd252788304, 'd263836680192, 'd15255162880, - 'd9694081024, 'd348975392, 'd269685833728, 'd8142476288, - 'd9587174400, 'd439889728, 'd271986458624, 'd1074818560, - 'd9375527936, 'd524595744, 'd270781579264, - 'd5866192896, - 'd9063308288, 'd602243328, 'd266154344448, - 'd12601840640, - 'd8655766528, 'd672076160, 'd258226323456, - 'd19057170432, - 'd8159164928, 'd733439296, 'd247155507200, - 'd25161789440, - 'd7580680704, 'd785784512, 'd233133752320, - 'd30850611200, - 'd6928315392, 'd828675456, 'd216383995904, - 'd36064505856, - 'd6210783744, 'd861790464, 'd197157126144, - 'd40750891008, - 'd5437403136, 'd884924608, 'd175728607232, - 'd44864233472, - 'd4617976320, 'd897990272, 'd152394776576, - 'd48366440448, - 'd3762670080, 'd901015872, 'd127469125632, - 'd51227189248, - 'd2881891584, 'd894144000, 'd101278294016, - 'd53424144384, - 'd1986164096, 'd877627648, 'd74158080000, - 'd54943068160, - 'd1086004096, 'd851825792, 'd46449369088, - 'd55777853440, - 'd191799792, 'd817197120, 'd18494062592, - 'd55930470400, 'd686306496, 'd774293504, - 'd9368892416, - 'd55410786304, 'd1538531200, 'd723751744, - 'd36807413760, - 'd54236319744, 'd2355556864, 'd666285184, - 'd63500029952, - 'd52431921152, 'd3128631040, 'd602673856, - 'd89139437568, - 'd50029350912, 'd3849658368, 'd533754816, - 'd113435836416, - 'd47066787840, 'd4511283200, 'd460411168, - 'd136120008704, - 'd43588292608, 'd5106960896, 'd383561312, - 'd156946137088, - 'd39643185152, 'd5631021568, 'd304147840, - 'd175694184448, - 'd35285385216, 'd6078718976, 'd223126112, - 'd192172146688, - 'd30572709888, 'd6446269952, 'd141453168, - 'd206217691136, - 'd25566150656, 'd6730883584, 'd60076656, - 'd217699647488, - 'd20329084928, 'd6930774016, - 'd20075964, - 'd226518974464, - 'd14926526464, 'd7045166592, - 'd98107728, - 'd232609366016, - 'd9424327680, 'd7074288128, - 'd173161984, - 'd235937497088, - 'd3888407296, 'd7019345920, - 'd244431584, - 'd236502859776, 'd1616015232, 'd6882502144, - 'd311167360, - 'd234337206272, 'd7025165824, 'd6666826240, - 'd372685728, - 'd229503696896, 'd12277432320, 'd6376248320, - 'd428375552, - 'd222095589376, 'd17314041856, 'd6015498752, - 'd477703744, - 'd212234715136, 'd22079696896, 'd5590036992, - 'd520220320, - 'd200069513216, 'd26523152384, 'd5105980416, - 'd555562048, - 'd185772982272, 'd30597754880, 'd4570017280, - 'd583455104, - 'd169540141056, 'd34261897216, 'd3989324800, - 'd603716864, - 'd151585505280, 'd37479415808, 'd3371473408, - 'd616256256, - 'd132140228608, 'd40219930624, 'd2724335104, - 'd621073344, - 'd111449161728, 'd42459090944, 'd2055986048, - 'd618257728, - 'd89767772160, 'd44178755584, 'd1374610176, - 'd607985920, - 'd67359031296, 'd45367111680, 'd688401792, - 'd590518080, - 'd44490215424, 'd46018699264, 'd5471468, - 'd566193024, - 'd21429762048, 'd46134370304, - 'd666247424, - 'd535423520, 'd1555883136, 'd45721169920, - 'd1319086976, - 'd498689888, 'd24205301760, 'd44792164352, - 'd1945729536, - 'd456533408, 'd46265061376, 'd43366166528, - 'd2539286272, - 'd409548928, 'd67492519936, 'd41467457536, - 'd3093369600, - 'd358377120, 'd87658446848, 'd39125377024, - 'd3602159872, - 'd303696256, 'd106549485568, 'd36373929984, - 'd4060461568, - 'd246213632, 'd123970330624, 'd33251299328, - 'd4463754240, - 'd186656976, 'd139745705984, 'd29799337984, - 'd4808232448, - 'd125765560, 'd153722093568, 'd26063024128, - 'd5090839552, - 'd64281496, 'd165769084928, 'd22089889792, - 'd5309289472, - 'd2941044, 'd175780577280, 'd17929424896, - 'd5462078464, 'd57533836, 'd183675584512, 'd13632480256, - 'd5548493312, 'd116443600, 'd189398745088, 'd9250644992, - 'd5568603136, 'd173118880, 'd192920535040, 'd4835645952, - 'd5523246592, 'd226927712, 'd194237251584, 'd438742560, - 'd5414009344, 'd277282272, 'd193370537984, - 'd3889856000, - 'd5243192832, 'd323644960, 'd190366760960, - 'd8101555712, - 'd5013775360, 'd365533728, 'd185296093184, - 'd12149912576, - 'd4729367040, 'd402526848, 'd178251268096, - 'd15991135232, - 'd4394157056, 'd434266688, 'd169346187264, - 'd19584544768, - 'd4012854528, 'd460462816, 'd158714167296, - 'd22892994560, - 'd3590626816, 'd480894272, 'd146506186752, - 'd25883242496, - 'd3133030656, 'd495411008, 'd132888772608, - 'd28526272512, - 'd2645941760, 'd503934304, 'd118041862144, - 'd30797553664, - 'd2135481216, 'd506456576, 'd102156492800, - 'd32677253120, - 'd1607940736, 'd503040352, 'd85432393728, - 'd34150387712, - 'd1069706688, 'd493816192, 'd68075581440, - 'd35206914048, - 'd527184576, 'd478980192, 'd50295820288, - 'd35841761280, 'd13275691, 'd458790528, 'd32304191488, - 'd36054810624, 'd545452224, 'd433563520, 'd14310600704, - 'd35850821632, 'd1063321216, 'd403668896, - 'd3478606336, - 'd35239272448, 'd1561123456, 'd369524608, - 'd20862973952, - 'd34234189824, 'd2033426688, 'd331591296, - 'd37650149376, - 'd32853913600, 'd2475182848, 'd290366144, - 'd53657956352, - 'd31120795648, 'd2881780480, 'd246376544, - 'd68716351488, - 'd29060892672, 'd3249091072, 'd200173424, - 'd82669150208, - 'd26703589376, 'd3573507840, 'd152324528, - 'd95375622144, - 'd24081211392, 'd3851980032, 'd103407576, - 'd106711851008, - 'd21228597248, 'd4082038528, 'd54003312, - 'd116571865088, - 'd18182653952, 'd4261814272, 'd4688806, - 'd124868567040, - 'd14981902336, 'd4390051328, - 'd43969216, - 'd131534446592, - 'd11665993728, 'd4466109440, - 'd91420760, - 'd136521965568, - 'd8275239936, 'd4489962496, - 'd137138640, - 'd139803836416, - 'd4850135552, 'd4462188544, - 'd180624272, - 'd141372964864, - 'd1430882688, 'd4383951872, - 'd221412864, - 'd141242171392, 'd1943064960, 'd4256981760, - 'd259078384, - 'd139443732480, 'd5233448448, 'd4083541248, - 'd293237696, - 'd136028684288, 'd8403623936, 'd3866393344, - 'd323554464, - 'd131065856000, 'd11418961920, 'd3608760064, - 'd349742080, - 'd124640845824, 'd14247211008, 'd3314277632, - 'd371566368, - 'd116854710272, 'd16858833920, 'd2986947328, - 'd388847200, - 'd107822514176, 'd19227299840, 'd2631084288, - 'd401459936, - 'd97671798784, 'd21329344512, 'd2251260672, - 'd409335712, - 'd86540869632, 'd23145181184, 'd1852249216, - 'd412461504, - 'd74577018880, 'd24658677760, 'd1438965504, - 'd410879232, - 'd61934665728, 'd25857468416, 'd1016407424, - 'd404684448, - 'd48773451776, 'd26733047808, 'd589596736, - 'd394024256, - 'd35256303616, 'd27280797696, 'd163520480, - 'd379094880, - 'd21547479040, 'd27499972608, - 'd256926192, - 'd360138432, - 'd7810651136, 'd27393648640, - 'd666995136, - 'd337439520, 'd5792974336, 'd26968619008, - 'd1062137472, - 'd311321088, 'd19106494464, 'd26235260928, - 'd1438052992, - 'd282140192, 'd31979048960, 'd25207339008, - 'd1790736000, - 'd250283168, 'd44267466752, 'd23901808640, - 'd2116516096, - 'd216160832, 'd55837798400, 'd22338547712, - 'd2412095488, - 'd180203184, 'd66566709248, 'd20540094464, - 'd2674580480, - 'd142854208, 'd76342730752, 'd18531325952, - 'd2901509120, - 'd104566496, 'd85067358208, 'd16339141632, - 'd3090871296, - 'd65795828, 'd92655960064, 'd13992113152, - 'd3241124864, - 'd26995910, 'd99038543872, 'd11520123904, - 'd3351205888, 'd11386859, 'd104160296960, 'd8954007552, - 'd3420532224, 'd48918428, 'd107981996032, 'd6325167616, - 'd3449003264, 'd85181896, 'd110480179200, 'd3665207808, - 'd3436992256, 'd119782032, 'd111647170560, 'd1005561408, - 'd3385333760, 'd152349504, 'd111490867200, - 'd1622868352, - 'd3295307008, 'd182544688, 'd110034436096, - 'd4190059008, - 'd3168613632, 'd210061120, 'd107315757056, - 'd6667201024, - 'd3007350016, 'd234628432, 'd103386734592, - 'd9027011584, - 'd2813977088, 'd256014944, 'd98312503296, - 'd11244024832, - 'd2591285760, 'd274029632, 'd92170379264, - 'd13294855168, - 'd2342358784, 'd288523648, 'd85048827904, - 'd15158435840, - 'd2070530560, 'd299391392, 'd77046226944, - 'd16816222208, - 'd1779343616, 'd306570976, 'd68269547520, - 'd18252363776, - 'd1472505088, 'd310044160, 'd58832982016, - 'd19453847552, - 'd1153840384, 'd309835904, 'd48856506368, - 'd20410593280, - 'd827246976, 'd306013216, 'd38464389120, - 'd21115523072, - 'd496648352, 'd298683904, 'd27783663616, - 'd21564604416, - 'd165947968, 'd287994368, 'd16942639104, - 'd21756829696, 'd161015488, 'd274127456, 'd6069367296, - 'd21694183424, 'd480511552, 'd257299680, - 'd4709823488, - 'd21381576704, 'd788959168, 'd237758064, - 'd15271768064, - 'd20826730496, 'd1082965888, 'd215776896, - 'd25497839616, - 'd20040044544, 'd1359363712, 'd191653968, - 'd35275247616, - 'd19034429440, 'd1615242112, 'd165706880, - 'd44498239488, - 'd17825124352, 'd1847977472, 'd138268864, - 'd53069225984, - 'd16429464576, 'd2055258368, 'd109684824, - 'd60899762176, - 'd14866663424, 'd2235107584, 'd80307000, - 'd67911417856, - 'd13157547008, 'd2385898752, 'd50490892, - 'd74036527104, - 'd11324291072, 'd2506369792, 'd20591002, - 'd79218802688, - 'd9390139392, 'd2595631104, - 'd9043209, - 'd83413778432, - 'd7379118592, 'd2653169920, - 'd38071296, - 'd86589120512, - 'd5315746304, 'd2678849792, - 'd66165620, - 'd88724840448, - 'd3224739072, 'd2672905216, - 'd93014920, - 'd89813286912, - 'd1130721792, 'd2635934208, - 'd118327656, - 'd89859039232, 'd942053824, 'd2568883456, - 'd141835040, - 'd88878645248, 'd2969985280, 'd2473032960, - 'd163293760, - 'd86900252672, 'd4930381312, 'd2349974784, - 'd182488384, - 'd83963068416, 'd6801708544, 'd2201590016, - 'd199233408, - 'd80116711424, 'd8563822592, 'd2030020992, - 'd213374832, - 'd75420508160, 'd10198177792, 'd1837643904, - 'd224791472, - 'd69942599680, 'd11688014848, 'd1627035520, - 'd233395808, - 'd63759036416, 'd13018524672, 'd1400941312, - 'd239134400, - 'd56952745984, 'd14176988160, 'd1162240128, - 'd241988000, - 'd49612476416, 'd15152887808, 'd913908864, - 'd241971088, - 'd41831669760, 'd15937992704, 'd658986304, - 'd239131280, - 'd33707284480, 'd16526415872, 'd400536864, - 'd233548080, - 'd25338644480, 'd16914642944, 'd141614768, - 'd225331520, - 'd16826230784, 'd17101535232, - 'd114771248, - 'd214620368, - 'd8270504960, 'd17088299008, - 'd365691968, - 'd201579968, 'd229250672, 'd16878435328, - 'd608330368, - 'd186399968, 'd8576060928, 'd16477662208, - 'd840012160, - 'd169291648, 'd16676343808, 'd15893807104, - 'd1058234624, - 'd150485136, 'd24440932352, 'd15136688128, - 'd1260692480, - 'd130226448, 'd31786033152, 'd14217958400, - 'd1445301760, - 'd108774312, 'd38634110976, 'd13150946304, - 'd1610219392, - 'd86397032, 'd44914671616, 'd11950475264, - 'd1753861248, - 'd63369172, 'd50564964352, 'd10632657920, - 'd1874915968, - 'd39968276, 'd55530573824, 'd9214700544, - 'd1972355584, - 'd16471616, 'd59765919744, 'd7714673664, - 'd2045442560, 'd6847026, 'd63234625536, 'd6151298560, - 'd2093733376, 'd29720462, 'd65909788672, 'd4543711744, - 'd2117079296, 'd51891092, 'd67774132224, 'd2911243008, - 'd2115622528, 'd73113720, 'd68820041728, 'd1273183616, - 'd2089790208, 'd93158192, 'd69049499648, - 'd351433280, - 'd2040284416, 'd111811808, 'd68473896960, - 'd1944049536, - 'd1968069376, 'd128881496, 'd67113725952, - 'd3486789120, - 'd1874356352, 'd144195728, 'd64998219776, - 'd4962652672, - 'd1760584960, 'd157606112, 'd62164844544, - 'd6355700736, - 'd1628403200, 'd168988784, 'd58658750464, - 'd7651218944, - 'd1479644416, 'd178245392, 'd54532087808, - 'd8835868672, - 'd1316303360, 'd185303792, 'd49843318784, - 'd9897820160, - 'd1140510208, 'd190118496, 'd44656418816, - 'd10826858496, - 'd954503680, 'd192670752, 'd39040032768, - 'd11614480384, - 'd760603392, 'd192968256, 'd33066635264, - 'd12253963264, - 'd561181504, 'd191044672, 'd26811590656, - 'd12740410368, - 'd358634592, 'd186958800, 'd20352258048, - 'd13070778368, - 'd155355344, 'd180793488, 'd13767048192, - 'd13243881472, 'd46295076, 'd172654240, 'd7134508032, - 'd13260374016, 'd244013680, 'd162667648, 'd532402080, - 'd13122712576, 'd435581472, 'd150979568, - 'd5963171840, - 'd12835095552, 'd618887680, 'd137753088, - 'd12278635520, - 'd12403388416, 'd791952384, 'd123166384, - 'd18343737344, - 'd11835023360, 'd952947136, 'd107410400, - 'd24092315648, - 'd11138892800, 'd1100213760, 'd90686408, - 'd29462990848, - 'd10325217280, 'd1232280576, 'd73203528, - 'd34399793152, - 'd9405405184, 'd1347876480, 'd55176152, - 'd38852730880, - 'd8391904768, 'd1445942016, 'd36821416, - 'd42778251264, - 'd7298036736, 'd1525638272, 'd18356602, - 'd46139658240, - 'd6137830912, 'd1586352896, - 'd3364, - 'd48907403264, - 'd4925849088, 'd1627703296, - 'd18048354, - 'd51059314688, - 'd3677007104, 'd1649537408, - 'd35575396, - 'd52580737024, - 'd2406398464, 'd1651931392, - 'd52390896, - 'd53464559616, - 'd1129114624, 'd1635185152, - 'd68312728, - 'd53711183872, 'd139928944, 'd1599814784, - 'd83172152, - 'd53328396288, 'd1386162304, 'd1546543488, - 'd96815528, - 'd52331134976, 'd2595524096, 'd1476289152, - 'd109105848, - 'd50741219328, 'd3754616064, 'd1390150784, - 'd119924056, - 'd48586973184, 'd4850846208, 'd1289392896, - 'd129170104, - 'd45902774272, 'd5872562688, 'd1175427840, - 'd136763808, - 'd42728583168, 'd6809170432, 'd1049796992, - 'd142645424, - 'd39109353472, 'd7651239424, 'd914150976, - 'd146776032, - 'd35094458368, 'd8390590464, 'd770228544, - 'd149137584, - 'd30737025024, 'd9020372992, 'd619834944, - 'd149732832, - 'd26093264896, 'd9535118336, 'd464820192, - 'd148584864, - 'd21221765120, 'd9930782720, 'd307056544, - 'd145736576, - 'd16182777856, 'd10204768256, 'd148416656, - 'd141249808, - 'd11037487104, 'd10355931136, - 'd9248055, - 'd135204288, - 'd5847291392, 'd10384567296, - 'd164128624, - 'd127696448, - 'd673083584, 'd10292387840, - 'd314478656, - 'd118838032, 'd4425443328, 'd10082473984, - 'd458633504, - 'd108754496, 'd9390467072, 'd9759219712, - 'd595028224, - 'd97583376, 'd14166675456, 'd9328256000, - 'd722214016, - 'd85472480, 'd18701864960, 'd8796367872, - 'd838872960, - 'd72578000, 'd22947489792, 'd8171397632, - 'd943831040, - 'd59062548, 'd26859171840, 'd7462130688, - 'd1036069504, - 'd45093212, 'd30397132800, 'd6678184448, - 'd1114734080, - 'd30839494, 'd33526589440, 'd5829879808, - 'd1179141760, - 'd16471352, 'd36218060800, 'd4928109056, - 'd1228786048, - 'd2157196, 'd38447636480, 'd3984203008, - 'd1263340160, 'd11938022, 'd40197140480, 'd3009790464, - 'd1282657280, 'd25654662, 'd41454268416, 'd2016659712, - 'd1286769408, 'd38840152, 'd42212614144, 'd1016618176, - 'd1275884288, 'd51350640, 'd42471653376, 'd21356334, - 'd1250379776, 'd63052516, 'd42236645376, - 'd957685888, - 'd1210796416, 'd73823768, 'd41518489600, - 'd1909447296, - 'd1157828864, 'd83555224, 'd40333484032, - 'd2823367424, - 'd1092315392, 'd92151592, 'd38703067136, - 'd3689500160, - 'd1015224960, 'd99532312, 'd36653469696, - 'd4498618368, - 'd927644736, 'd105632264, 'd34215340032, - 'd5242309120, - 'd830765056, 'd110402272, 'd31423309824, - 'd5913057792, - 'd725863872, 'd113809368, 'd28315527168, - 'd6504319488, - 'd614290688, 'd115836928, 'd24933158912, - 'd7010576896, - 'd497449664, 'd116484592, 'd21319860224, - 'd7427391488, - 'd376782464, 'd115767992, 'd17521235968, - 'd7751432704, - 'd253750912, 'd113718288, 'd13584269312, - 'd7980498432, - 'd129819680, 'd110381560, 'd9556759552, - 'd8113524224, - 'd6439408, 'd105818040, 'd5486758400, - 'd8150574080, 'd114969968, 'd100101136, 'd1422006400, - 'd8092821504, 'd233035072, 'd93316416, - 'd2590614528, - 'd7942518272, 'd346444256, 'd85560352, - 'd6505608704, - 'd7702948864, 'd453961664, 'd76939064, - 'd10279368704, - 'd7378376192, 'd554440448, 'd67566928, - 'd13870651392, - 'd6973975552, 'd646834304, 'd57565096, - 'd17241012224, - 'd6495759872, 'd730208128, 'd47059976, - 'd20355205120, - 'd5950494720, 'd803746816, 'd36181704, - 'd23181537280, - 'd5345609216, 'd866762944, 'd25062552, - 'd25692176384, - 'd4689098240, 'd918702144, 'd13835381, - 'd27863408640, - 'd3989420544, 'd959147840, 'd2632072, - 'd29675841536, - 'd3255392000, 'd987823232, - 'd8417969, - 'd31114557440, - 'd2496078848, 'd1004592512, - 'd19189274, - 'd32169211904, - 'd1720688896, 'd1009460096, - 'd29561700, - 'd32834078720, - 'd938460864, 'd1002568000, - 'd39421732, - 'd33108035584, - 'd158558640, 'd984192000, - 'd48663680, - 'd32994498560, 'd610034432, 'd954736192, - 'd57190776};
	localparam logic signed[63:0] hb[0:1999] = {'d7033096503296, 'd32897980416, - 'd10967230464, - 'd63928604, 'd7000245665792, 'd98394423296, - 'd10337267712, - 'd188110032, 'd6934845456384, 'd162997501952, - 'd9086782464, - 'd301512896, 'd6837488844800, 'd226124627968, - 'd7233756672, - 'd397524544, 'd6709056110592, 'd287210536960, - 'd4804252672, - 'd470098240, 'd6550703833088, 'd345713672192, - 'd1831931776, - 'd513814560, 'd6363853881344, 'd401122131968, 'd1642511488, - 'd523933696, 'd6150172966912, 'd452959338496, 'd5571985920, - 'd496438560, 'd5911558488064, 'd500788854784, 'd9903706112, - 'd428068320, 'd5650113888256, 'd544219168768, 'd14579948544, - 'd316342016, 'd5368126111744, 'd582907527168, 'd19538849792, - 'd159572240, 'd5068042010624, 'd616563212288, 'd24715249664, 'd43130884, 'd4752438460416, 'd644950327296, 'd30041542656, 'd291865696, 'd4423997194240, 'd667889827840, 'd35448557568, 'd585954240, 'd4085474918400, 'd685260537856, 'd40866439168, 'd923966848, 'd3739673690112, 'd697000263680, 'd46225510400, 'd1303755136, 'd3389412343808, 'd703105531904, 'd51457126400, 'd1722493184, 'd3037497131008, 'd703630671872, 'd56494514176, 'd2176726784, 'd2686692360192, 'd698686832640, 'd61273546752, 'd2662427904, 'd2339693658112, 'd688439820288, 'd65733513216, 'd3175056896, 'd1999099920384, 'd673107279872, 'd69817778176, 'd3709628672, 'd1667389456384, 'd652956008448, 'd73474457600, 'd4260784384, 'd1346895216640, 'd628297957376, 'd76656959488, 'd4822863872, 'd1039784017920, 'd599486234624, 'd79324479488, 'd5389984768, 'd748036685824, 'd566910648320, 'd81442447360, 'd5956117504, 'd473431015424, 'd530992660480, 'd82982838272, 'd6515166720, 'd217527091200, 'd492180406272, 'd83924451328, 'd7061048320, - 'd18344486912, 'd450943287296, 'd84253073408, 'd7587765248, - 'd233092038656, 'd407766368256, 'd83961561088, 'd8089484800, - 'd425869180928, 'd363144806400, 'd83049857024, 'd8560607232, - 'd596078428160, 'd317578280960, 'd81524924416, 'd8995835904, - 'd743372095488, 'd271565209600, 'd79400542208, 'd9390236672, - 'd867650306048, 'd225597456384, 'd76697108480, 'd9739302912, - 'd969056190464, 'd180154810368, 'd73441320960, 'd10038998016, - 'd1047968874496, 'd135700045824, 'd69665783808, 'd10285808640, - 'd1104993583104, 'd92673966080, 'd65408569344, 'd10476781568, - 'd1140949254144, 'd51490967552, 'd60712722432, 'd10609551360, - 'd1156854972416, 'd12534914048, 'd55625695232, 'd10682369024, - 'd1153913061376, - 'd23844581376, 'd50198769664, 'd10694119424, - 'd1133491388416, - 'd57335398400, 'd44486422528, 'd10644324352, - 'd1097103966208, - 'd87665672192, 'd38545653760, 'd10533150720, - 'd1046390308864, - 'd114606071808, 'd32435316736, 'd10361399296, - 'd983093477376, - 'd137971515392, 'd26215440384, 'd10130492416, - 'd909037731840, - 'd157622370304, 'd19946518528, 'd9842454528, - 'd826105724928, - 'd173465124864, 'd13688829952, 'd9499883520, - 'd736215171072, - 'd185452544000, 'd7501764608, 'd9105917952, - 'd641296105472, - 'd193583169536, 'd1443165440, 'd8664196096, - 'd543267749888, - 'd197900484608, - 'd4431298048, 'd8178812416, - 'd444016885760, - 'd198491455488, - 'd10068722688, 'd7654265856, - 'd345376227328, - 'd195484614656, - 'd15419525120, 'd7095408640, - 'd249104269312, - 'd189047783424, - 'd20437946368, 'd6507388928, - 'd156866412544, - 'd179385237504, - 'd25082505216, 'd5895589888, - 'd70217392128, - 'd166734675968, - 'd29316399104, 'd5265568768, 'd9414508544, - 'd151363747840, - 'd33107843072, 'd4622995968, 'd80741564416, - 'd133566259200, - 'd36430344192, 'd3973589248, 'd142628683776, - 'd113658347520, - 'd39262916608, 'd3323052544, 'd194103558144, - 'd91974221824, - 'd41590218752, 'd2677014272, 'd234364616704, - 'd68861943808, - 'd43402641408, 'd2040966400, 'd262786842624, - 'd44679032832, - 'd44696309760, 'd1420208256, 'd278925475840, - 'd19788113920, - 'd45473042432, 'd819790720, 'd282517438464, 'd5447470592, - 'd45740224512, 'd244465792, 'd273480531968, 'd30667960320, - 'd45510623232, - 'd301360416, 'd251910750208, 'd55521345536, - 'd44802162688, - 'd813669824, 'd218077265920, 'd79667380224, - 'd43637624832, - 'd1288869760, 'd172415664128, 'd102781378560, - 'd42044309504, - 'd1723824640, 'd115519225856, 'd124557795328, - 'd40053633024, - 'd2115882240, 'd48128520192, 'd144713433088, - 'd37700722688, - 'd2462894336, - 'd28880474112, 'd162990424064, - 'd35023921152, - 'd2763230464, - 'd114509742080, 'd179158859776, - 'd32064319488, - 'd3015787008, - 'd207653748736, 'd193018920960, - 'd28865234944, - 'd3219988736, - 'd307115032576, 'd204402835456, - 'd25471664128, - 'd3375784960, - 'd411620442112, 'd213176172544, - 'd21929756672, - 'd3483641344, - 'd519838269440, 'd219238973440, - 'd18286260224, - 'd3544522240, - 'd630395568128, 'd222526259200, - 'd14587981824, - 'd3559872512, - 'd741895634944, 'd223008227328, - 'd10881244160, - 'd3531590144, - 'd852935704576, 'd220690022400, - 'd7211374080, - 'd3461996544, - 'd962124054528, 'd215611097088, - 'd3622200320, - 'd3353801728, - 'd1068097273856, 'd207844130816, - 'd155578656, - 'd3210066176, - 'd1169536057344, 'd197493669888, 'd3149049344, - 'd3034159104, - 'd1265181130752, 'd184694308864, 'd6255063040, - 'd2829713920, - 'd1353847668736, 'd169608675328, 'd9129030656, - 'd2600581376, - 'd1434438467584, 'd152425005056, 'd11741032448, - 'd2350781696, - 'd1505956593664, 'd133354577920, 'd14064936960, - 'd2084455552, - 'd1567515475968, 'd112628752384, 'd16078633984, - 'd1805813376, - 'd1618349129728, 'd90496016384, 'd17764208640, - 'd1519086592, - 'd1657819234304, 'd67218747392, 'd19108071424, - 'd1228478592, - 'd1685421162496, 'd43069902848, 'd20101029888, - 'd938116672, - 'd1700789092352, 'd18329671680, 'd20738314240, - 'd652006464, - 'd1703698104320, - 'd6717959680, 'd21019545600, - 'd373988160, - 'd1694065885184, - 'd31788576768, 'd20948656128, - 'd107695488, - 'd1671951417344, - 'd56600698880, 'd20533766144, 'd143481952, - 'd1637553012736, - 'd80879017984, 'd19787003904, 'd376432992, - 'd1591204642816, - 'd104357543936, 'd18724286464, 'd588355264, - 'd1533370171392, - 'd126782562304, 'd17365071872, 'd776781440, - 'd1464636669952, - 'd147915423744, 'd15732052992, 'd939601280, - 'd1385706160128, - 'd167535099904, 'd13850836992, 'd1075078784, - 'd1297386569728, - 'd185440518144, 'd11749591040, 'd1181864704, - 'd1200580722688, - 'd201452535808, 'd9458661376, 'd1259004928, - 'd1096275197952, - 'd215415816192, 'd7010174464, 'd1305943424, - 'd985527877632, - 'd227200188416, 'd4437632000, 'd1322520576, - 'd869455364096, - 'd236701794304, 'd1775485824, 'd1308967168, - 'd749219348480, - 'd243843940352, - 'd941283776, 'd1265894400, - 'd626012913664, - 'd248577572864, - 'd3677590016, 'd1194278144, - 'd501046935552, - 'd250881425408, - 'd6398656512, 'd1095440768, - 'd375535730688, - 'd250761838592, - 'd9070423040, 'd971028672, - 'd250683834368, - 'd248252301312, - 'd11659934720, 'd822986240, - 'd127672295424, - 'd243412647936, - 'd14135713792, 'd653526912, - 'd7645917696, - 'd236328009728, - 'd16468104192, 'd465101920, 'd108299083776, - 'd227107389440, - 'd18629595136, 'd260366176, 'd219126661120, - 'd215882104832, - 'd20595109888, 'd42143052, 'd323871637504, - 'd202803920896, - 'd22342254592, - 'd186612704, 'd421649350656, - 'd188043018240, - 'd23851552768, - 'd422852640, 'd511664455680, - 'd171785748480, - 'd25106614272, - 'd663472896, 'd593218240512, - 'd154232242176, - 'd26094284800, - 'd905352320, 'd665715081216, - 'd135593918464, - 'd26804754432, - 'd1145390336, 'd728667193344, - 'd116090904576, - 'd27231608832, - 'd1380543744, 'd781698727936, - 'd95949373440, - 'd27371864064, - 'd1607862400, 'd824547606528, - 'd75398856704, - 'd27225939968, - 'd1824522752, 'd857067028480, - 'd54669598720, - 'd26797602816, - 'd2027859968, 'd879224750080, - 'd33989888000, - 'd26093875200, - 'd2215397376, 'd891101773824, - 'd13583513600, - 'd25124898816, - 'd2384873216, 'd892889333760, 'd6332733440, - 'd23903772672, - 'd2534263552, 'd884884701184, 'd25551407104, - 'd22446352384, - 'd2661804288, 'd867486269440, 'd43876618240, - 'd20771020800, - 'd2766007296, 'd841186934784, 'd61126078464, - 'd18898444288, - 'd2845674240, 'd806566887424, 'd77132947456, - 'd16851289088, - 'd2899907328, 'd764285681664, 'd91747483648, - 'd14653930496, - 'd2928114688, 'd715073060864, 'd104838455296, - 'd12332148736, - 'd2930013696, 'd659719585792, 'd116294311936, - 'd9912799232, - 'd2905629696, 'd599066345472, 'd126024146944, - 'd7423496704, - 'd2855291904, 'd533994668032, 'd133958361088, - 'd4892274176, - 'd2779624704, 'd465415241728, 'd140049088512, - 'd2347257600, - 'd2679536640, 'd394257203200, 'd144270393344, 'd183660272, - 'd2556206336, 'd321457225728, 'd146618138624, 'd2673139712, - 'd2411064576, 'd247948623872, 'd147109675008, 'd5094700032, - 'd2245774336, 'd174650785792, 'd145783259136, 'd7423012352, - 'd2062207744, 'd102458908672, 'd142697250816, 'd9634170880, - 'd1862423296, 'd32234213376, 'd137929080832, 'd11705949184, - 'd1648637312, - 'd35205341184, 'd131574038528, 'd13618027520, - 'd1423197824, - 'd99093577728, 'd123743797248, 'd15352196096, - 'd1188554880, - 'd158723964928, 'd114564939776, 'd16892532736, - 'd947231424, - 'd213456617472, 'd104177123328, 'd18225549312, - 'd701792896, - 'd262724354048, 'd92731334656, 'd19340306432, - 'd454817568, - 'd306037915648, 'd80387866624, 'd20228497408, - 'd208866800, - 'd342990127104, 'd67314339840, 'd20884506624, 'd33544018, - 'd373259010048, 'd53683642368, 'd21305427968, 'd269973504, - 'd396609880064, 'd39671808000, 'd21491048448, 'd498081024, - 'd412896460800, 'd25455941632, 'd21443817472, 'd715651776, - 'd422060851200, 'd11212149760, 'd21168769024, 'd920620160, - 'd424132542464, - 'd2886491648, 'd20673421312, 'd1111091072, - 'd419226353664, - 'd16671883264, 'd19967651840, 'd1285358592, - 'd407539548160, - 'd29982767104, 'd19063545856, 'd1441922816, - 'd389347966976, - 'd42666471424, 'd17975222272, 'd1579503232, - 'd365001244672, - 'd54580543488, 'd16718628864, 'd1697049984, - 'd334917435392, - 'd65594208256, 'd15311344640, 'd1793752448, - 'd299576754176, - 'd75589697536, 'd13772339200, 'd1869043840, - 'd259514777600, - 'd84463378432, 'd12121732096, 'd1922604416, - 'd215315218432, - 'd92126724096, 'd10380551168, 'd1954360704, - 'd167602061312, - 'd98507071488, 'd8570467840, 'd1964482176, - 'd117031575552, - 'd103548190720, 'd6713540096, 'd1953375744, - 'd64283930624, - 'd107210645504, 'd4831954432, 'd1921676416, - 'd10054776832, - 'd109471981568, 'd2947766016, 'd1870237312, 'd44953247744, - 'd110326685696, 'd1082651264, 'd1800114816, 'd100038934528, - 'd109785948160, - 'd742337920, 'd1712554752, 'd154510770176, - 'd107877253120, - 'd2507003392, 'd1608973312, 'd207694921728, - 'd104643788800, - 'd4192218624, 'd1490939392, 'd258942943232, - 'd100143644672, - 'd5780130304, 'd1360152832, 'd307638960128, - 'd94448910336, - 'd7254341120, 'd1218423808, 'd353206403072, - 'd87644585984, - 'd8600073216, 'd1067649472, 'd395114184704, - 'd79827378176, - 'd9804311552, 'd909791232, 'd432882253824, - 'd71104356352, - 'd10855919616, 'd746850816, 'd466086363136, - 'd61591547904, - 'd11745739776, 'd580847104, 'd494362230784, - 'd51412426752, - 'd12466658304, 'd413792224, 'd517408784384, - 'd40696356864, - 'd13013656576, 'd247669072, 'd534990848000, - 'd29576974336, - 'd13383830528, 'd84408840, 'd546940780544, - 'd18190557184, - 'd13576387584, - 'd74130096, 'd553159360512, - 'd6674405888, - 'd13592614912, - 'd226182256, 'd553615949824, 'd4834780672, - 'd13435834368, - 'd370093632, 'd548347740160, 'd16202491904, - 'd13111324672, - 'd504338656, 'd537458442240, 'd27297931264, - 'd12626223104, - 'd627535488, 'd521115828224, 'd37995479040, - 'd11989416960, - 'd738459264, 'd499548880896, 'd48176078848, - 'd11211404288, - 'd836053504, 'd473044221952, 'd57728499712, - 'd10304146432, - 'd919438912, 'd441941950464, 'd66550517760, - 'd9280902144, - 'd987920768, 'd406630694912, 'd74549952512, - 'd8156052992, - 'd1040993088, 'd367542566912, 'd81645584384, - 'd6944914944, - 'd1078341504, 'd325147328512, 'd87767891968, - 'd5663543808, - 'd1099843200, 'd279946461184, 'd92859727872, - 'd4328539136, - 'd1105564672, 'd232466825216, 'd96876699648, - 'd2956838144, - 'd1095757824, 'd183254220800, 'd99787579392, - 'd1565513600, - 'd1070853440, 'd132866760704, 'd101574352896, - 'd171574784, - 'd1031453312, 'd81868210176, 'd102232301568, 'd1208231424, - 'd978319616, 'd30821447680, 'd101769781248, 'd2557609472, - 'd912363520, - 'd19718068224, 'd100207943680, 'd3860898560, - 'd834631680, - 'd69208547328, 'd97580294144, 'd5103242240, - 'd746291840, - 'd117127929856, 'd93932068864, 'd6270749696, - 'd648616768, - 'd162979545088, 'd89319563264, 'd7350639104, - 'd542967744, - 'd206297481216, 'd83809280000, 'd8331369472, - 'd430777056, - 'd246651437056, 'd77476986880, 'd9202753536, - 'd313529888, - 'd283651080192, 'd70406725632, 'd9956050944, - 'd192746128, - 'd316949954560, 'd62689660928, 'd10584052736, - 'd69961976, - 'd346248708096, 'd54422949888, 'd11081128960, 'd53288364, - 'd371297878016, 'd45708509184, 'd11443279872, 'd175490560, - 'd391899774976, 'd36651757568, 'd11668144128, 'd295167552, - 'd407910121472, 'd27360344064, 'd11755006976, 'd410896192, - 'd419238739968, 'd17942872064, 'd11704777728, 'd521323040, - 'd425849716736, 'd8507630592, 'd11519951872, 'd625179008, - 'd427760877568, - 'd838650880, 'd11204558848, 'd721292672, - 'd425042903040, - 'd9992007680, 'd10764085248, 'd808602688, - 'd417817427968, - 'd18852395008, 'd10205391872, 'd886167872, - 'd406254944256, - 'd27324768256, 'd9536608256, 'd953176704, - 'd390571982848, - 'd35320111104, 'd8767017984, 'd1008954368, - 'd371027836928, - 'd42756349952, 'd7906931200, 'd1052968640, - 'd347921055744, - 'd49559191552, 'd6967550976, 'd1084833536, - 'd321585086464, - 'd55662837760, 'd5960825344, 'd1104311424, - 'd292384145408, - 'd61010624512, 'd4899297280, 'd1111313664, - 'd260708253696, - 'd65555509248, 'd3795950592, 'd1105899136, - 'd226968616960, - 'd69260451840, 'd2664050688, 'd1088270976, - 'd191592300544, - 'd72098676736, 'd1516986752, 'd1058772032, - 'd155017199616, - 'd74053804032, 'd368114528, 'd1017878592, - 'd117686788096, - 'd75119886336, - 'd769398208, 'd966192896, - 'd80044908544, - 'd75301273600, - 'd1882721152, 'd904433792, - 'd42530721792, - 'd74612400128, - 'd2959504384, 'd833426688, - 'd5573702144, - 'd73077473280, - 'd3988013824, 'd754092160, 'd30411114496, - 'd70729965568, - 'd4957257216, 'd667433984, 'd65027657728, - 'd67612160000, - 'd5857098752, 'd574525888, 'd97903050752, - 'd63774429184, - 'd6678363136, 'd476498048, 'd128691486720, - 'd59274575872, - 'd7412924928, 'd374523168, 'd157077749760, - 'd54177009664, - 'd8053787136, 'd269802144, 'd182780313600, - 'd48551907328, - 'd8595142656, 'd163549664, 'd205553975296, - 'd42474287104, - 'd9032420352, 'd56980000, 'd225192067072, - 'd36023083008, - 'd9362321408, - 'd48707084, 'd241528176640, - 'd29280149504, - 'd9582834688, - 'd152339968, 'd254437326848, - 'd22329272320, - 'd9693236224, - 'd252788304, 'd263836680192, - 'd15255162880, - 'd9694081024, - 'd348975392, 'd269685833728, - 'd8142476288, - 'd9587174400, - 'd439889728, 'd271986458624, - 'd1074818560, - 'd9375527936, - 'd524595744, 'd270781579264, 'd5866192896, - 'd9063308288, - 'd602243328, 'd266154344448, 'd12601840640, - 'd8655766528, - 'd672076160, 'd258226323456, 'd19057170432, - 'd8159164928, - 'd733439296, 'd247155507200, 'd25161789440, - 'd7580680704, - 'd785784512, 'd233133752320, 'd30850611200, - 'd6928315392, - 'd828675456, 'd216383995904, 'd36064505856, - 'd6210783744, - 'd861790464, 'd197157126144, 'd40750891008, - 'd5437403136, - 'd884924608, 'd175728607232, 'd44864233472, - 'd4617976320, - 'd897990272, 'd152394776576, 'd48366440448, - 'd3762670080, - 'd901015872, 'd127469125632, 'd51227189248, - 'd2881891584, - 'd894144000, 'd101278294016, 'd53424144384, - 'd1986164096, - 'd877627648, 'd74158080000, 'd54943068160, - 'd1086004096, - 'd851825792, 'd46449369088, 'd55777853440, - 'd191799792, - 'd817197120, 'd18494062592, 'd55930470400, 'd686306496, - 'd774293504, - 'd9368892416, 'd55410786304, 'd1538531200, - 'd723751744, - 'd36807413760, 'd54236319744, 'd2355556864, - 'd666285184, - 'd63500029952, 'd52431921152, 'd3128631040, - 'd602673856, - 'd89139437568, 'd50029350912, 'd3849658368, - 'd533754816, - 'd113435836416, 'd47066787840, 'd4511283200, - 'd460411168, - 'd136120008704, 'd43588292608, 'd5106960896, - 'd383561312, - 'd156946137088, 'd39643185152, 'd5631021568, - 'd304147840, - 'd175694184448, 'd35285385216, 'd6078718976, - 'd223126112, - 'd192172146688, 'd30572709888, 'd6446269952, - 'd141453168, - 'd206217691136, 'd25566150656, 'd6730883584, - 'd60076656, - 'd217699647488, 'd20329084928, 'd6930774016, 'd20075964, - 'd226518974464, 'd14926526464, 'd7045166592, 'd98107728, - 'd232609366016, 'd9424327680, 'd7074288128, 'd173161984, - 'd235937497088, 'd3888407296, 'd7019345920, 'd244431584, - 'd236502859776, - 'd1616015232, 'd6882502144, 'd311167360, - 'd234337206272, - 'd7025165824, 'd6666826240, 'd372685728, - 'd229503696896, - 'd12277432320, 'd6376248320, 'd428375552, - 'd222095589376, - 'd17314041856, 'd6015498752, 'd477703744, - 'd212234715136, - 'd22079696896, 'd5590036992, 'd520220320, - 'd200069513216, - 'd26523152384, 'd5105980416, 'd555562048, - 'd185772982272, - 'd30597754880, 'd4570017280, 'd583455104, - 'd169540141056, - 'd34261897216, 'd3989324800, 'd603716864, - 'd151585505280, - 'd37479415808, 'd3371473408, 'd616256256, - 'd132140228608, - 'd40219930624, 'd2724335104, 'd621073344, - 'd111449161728, - 'd42459090944, 'd2055986048, 'd618257728, - 'd89767772160, - 'd44178755584, 'd1374610176, 'd607985920, - 'd67359031296, - 'd45367111680, 'd688401792, 'd590518080, - 'd44490215424, - 'd46018699264, 'd5471468, 'd566193024, - 'd21429762048, - 'd46134370304, - 'd666247424, 'd535423520, 'd1555883136, - 'd45721169920, - 'd1319086976, 'd498689888, 'd24205301760, - 'd44792164352, - 'd1945729536, 'd456533408, 'd46265061376, - 'd43366166528, - 'd2539286272, 'd409548928, 'd67492519936, - 'd41467457536, - 'd3093369600, 'd358377120, 'd87658446848, - 'd39125377024, - 'd3602159872, 'd303696256, 'd106549485568, - 'd36373929984, - 'd4060461568, 'd246213632, 'd123970330624, - 'd33251299328, - 'd4463754240, 'd186656976, 'd139745705984, - 'd29799337984, - 'd4808232448, 'd125765560, 'd153722093568, - 'd26063024128, - 'd5090839552, 'd64281496, 'd165769084928, - 'd22089889792, - 'd5309289472, 'd2941044, 'd175780577280, - 'd17929424896, - 'd5462078464, - 'd57533836, 'd183675584512, - 'd13632480256, - 'd5548493312, - 'd116443600, 'd189398745088, - 'd9250644992, - 'd5568603136, - 'd173118880, 'd192920535040, - 'd4835645952, - 'd5523246592, - 'd226927712, 'd194237251584, - 'd438742560, - 'd5414009344, - 'd277282272, 'd193370537984, 'd3889856000, - 'd5243192832, - 'd323644960, 'd190366760960, 'd8101555712, - 'd5013775360, - 'd365533728, 'd185296093184, 'd12149912576, - 'd4729367040, - 'd402526848, 'd178251268096, 'd15991135232, - 'd4394157056, - 'd434266688, 'd169346187264, 'd19584544768, - 'd4012854528, - 'd460462816, 'd158714167296, 'd22892994560, - 'd3590626816, - 'd480894272, 'd146506186752, 'd25883242496, - 'd3133030656, - 'd495411008, 'd132888772608, 'd28526272512, - 'd2645941760, - 'd503934304, 'd118041862144, 'd30797553664, - 'd2135481216, - 'd506456576, 'd102156492800, 'd32677253120, - 'd1607940736, - 'd503040352, 'd85432393728, 'd34150387712, - 'd1069706688, - 'd493816192, 'd68075581440, 'd35206914048, - 'd527184576, - 'd478980192, 'd50295820288, 'd35841761280, 'd13275691, - 'd458790528, 'd32304191488, 'd36054810624, 'd545452224, - 'd433563520, 'd14310600704, 'd35850821632, 'd1063321216, - 'd403668896, - 'd3478606336, 'd35239272448, 'd1561123456, - 'd369524608, - 'd20862973952, 'd34234189824, 'd2033426688, - 'd331591296, - 'd37650149376, 'd32853913600, 'd2475182848, - 'd290366144, - 'd53657956352, 'd31120795648, 'd2881780480, - 'd246376544, - 'd68716351488, 'd29060892672, 'd3249091072, - 'd200173424, - 'd82669150208, 'd26703589376, 'd3573507840, - 'd152324528, - 'd95375622144, 'd24081211392, 'd3851980032, - 'd103407576, - 'd106711851008, 'd21228597248, 'd4082038528, - 'd54003312, - 'd116571865088, 'd18182653952, 'd4261814272, - 'd4688806, - 'd124868567040, 'd14981902336, 'd4390051328, 'd43969216, - 'd131534446592, 'd11665993728, 'd4466109440, 'd91420760, - 'd136521965568, 'd8275239936, 'd4489962496, 'd137138640, - 'd139803836416, 'd4850135552, 'd4462188544, 'd180624272, - 'd141372964864, 'd1430882688, 'd4383951872, 'd221412864, - 'd141242171392, - 'd1943064960, 'd4256981760, 'd259078384, - 'd139443732480, - 'd5233448448, 'd4083541248, 'd293237696, - 'd136028684288, - 'd8403623936, 'd3866393344, 'd323554464, - 'd131065856000, - 'd11418961920, 'd3608760064, 'd349742080, - 'd124640845824, - 'd14247211008, 'd3314277632, 'd371566368, - 'd116854710272, - 'd16858833920, 'd2986947328, 'd388847200, - 'd107822514176, - 'd19227299840, 'd2631084288, 'd401459936, - 'd97671798784, - 'd21329344512, 'd2251260672, 'd409335712, - 'd86540869632, - 'd23145181184, 'd1852249216, 'd412461504, - 'd74577018880, - 'd24658677760, 'd1438965504, 'd410879232, - 'd61934665728, - 'd25857468416, 'd1016407424, 'd404684448, - 'd48773451776, - 'd26733047808, 'd589596736, 'd394024256, - 'd35256303616, - 'd27280797696, 'd163520480, 'd379094880, - 'd21547479040, - 'd27499972608, - 'd256926192, 'd360138432, - 'd7810651136, - 'd27393648640, - 'd666995136, 'd337439520, 'd5792974336, - 'd26968619008, - 'd1062137472, 'd311321088, 'd19106494464, - 'd26235260928, - 'd1438052992, 'd282140192, 'd31979048960, - 'd25207339008, - 'd1790736000, 'd250283168, 'd44267466752, - 'd23901808640, - 'd2116516096, 'd216160832, 'd55837798400, - 'd22338547712, - 'd2412095488, 'd180203184, 'd66566709248, - 'd20540094464, - 'd2674580480, 'd142854208, 'd76342730752, - 'd18531325952, - 'd2901509120, 'd104566496, 'd85067358208, - 'd16339141632, - 'd3090871296, 'd65795828, 'd92655960064, - 'd13992113152, - 'd3241124864, 'd26995910, 'd99038543872, - 'd11520123904, - 'd3351205888, - 'd11386859, 'd104160296960, - 'd8954007552, - 'd3420532224, - 'd48918428, 'd107981996032, - 'd6325167616, - 'd3449003264, - 'd85181896, 'd110480179200, - 'd3665207808, - 'd3436992256, - 'd119782032, 'd111647170560, - 'd1005561408, - 'd3385333760, - 'd152349504, 'd111490867200, 'd1622868352, - 'd3295307008, - 'd182544688, 'd110034436096, 'd4190059008, - 'd3168613632, - 'd210061120, 'd107315757056, 'd6667201024, - 'd3007350016, - 'd234628432, 'd103386734592, 'd9027011584, - 'd2813977088, - 'd256014944, 'd98312503296, 'd11244024832, - 'd2591285760, - 'd274029632, 'd92170379264, 'd13294855168, - 'd2342358784, - 'd288523648, 'd85048827904, 'd15158435840, - 'd2070530560, - 'd299391392, 'd77046226944, 'd16816222208, - 'd1779343616, - 'd306570976, 'd68269547520, 'd18252363776, - 'd1472505088, - 'd310044160, 'd58832982016, 'd19453847552, - 'd1153840384, - 'd309835904, 'd48856506368, 'd20410593280, - 'd827246976, - 'd306013216, 'd38464389120, 'd21115523072, - 'd496648352, - 'd298683904, 'd27783663616, 'd21564604416, - 'd165947968, - 'd287994368, 'd16942639104, 'd21756829696, 'd161015488, - 'd274127456, 'd6069367296, 'd21694183424, 'd480511552, - 'd257299680, - 'd4709823488, 'd21381576704, 'd788959168, - 'd237758064, - 'd15271768064, 'd20826730496, 'd1082965888, - 'd215776896, - 'd25497839616, 'd20040044544, 'd1359363712, - 'd191653968, - 'd35275247616, 'd19034429440, 'd1615242112, - 'd165706880, - 'd44498239488, 'd17825124352, 'd1847977472, - 'd138268864, - 'd53069225984, 'd16429464576, 'd2055258368, - 'd109684824, - 'd60899762176, 'd14866663424, 'd2235107584, - 'd80307000, - 'd67911417856, 'd13157547008, 'd2385898752, - 'd50490892, - 'd74036527104, 'd11324291072, 'd2506369792, - 'd20591002, - 'd79218802688, 'd9390139392, 'd2595631104, 'd9043209, - 'd83413778432, 'd7379118592, 'd2653169920, 'd38071296, - 'd86589120512, 'd5315746304, 'd2678849792, 'd66165620, - 'd88724840448, 'd3224739072, 'd2672905216, 'd93014920, - 'd89813286912, 'd1130721792, 'd2635934208, 'd118327656, - 'd89859039232, - 'd942053824, 'd2568883456, 'd141835040, - 'd88878645248, - 'd2969985280, 'd2473032960, 'd163293760, - 'd86900252672, - 'd4930381312, 'd2349974784, 'd182488384, - 'd83963068416, - 'd6801708544, 'd2201590016, 'd199233408, - 'd80116711424, - 'd8563822592, 'd2030020992, 'd213374832, - 'd75420508160, - 'd10198177792, 'd1837643904, 'd224791472, - 'd69942599680, - 'd11688014848, 'd1627035520, 'd233395808, - 'd63759036416, - 'd13018524672, 'd1400941312, 'd239134400, - 'd56952745984, - 'd14176988160, 'd1162240128, 'd241988000, - 'd49612476416, - 'd15152887808, 'd913908864, 'd241971088, - 'd41831669760, - 'd15937992704, 'd658986304, 'd239131280, - 'd33707284480, - 'd16526415872, 'd400536864, 'd233548080, - 'd25338644480, - 'd16914642944, 'd141614768, 'd225331520, - 'd16826230784, - 'd17101535232, - 'd114771248, 'd214620368, - 'd8270504960, - 'd17088299008, - 'd365691968, 'd201579968, 'd229250672, - 'd16878435328, - 'd608330368, 'd186399968, 'd8576060928, - 'd16477662208, - 'd840012160, 'd169291648, 'd16676343808, - 'd15893807104, - 'd1058234624, 'd150485136, 'd24440932352, - 'd15136688128, - 'd1260692480, 'd130226448, 'd31786033152, - 'd14217958400, - 'd1445301760, 'd108774312, 'd38634110976, - 'd13150946304, - 'd1610219392, 'd86397032, 'd44914671616, - 'd11950475264, - 'd1753861248, 'd63369172, 'd50564964352, - 'd10632657920, - 'd1874915968, 'd39968276, 'd55530573824, - 'd9214700544, - 'd1972355584, 'd16471616, 'd59765919744, - 'd7714673664, - 'd2045442560, - 'd6847026, 'd63234625536, - 'd6151298560, - 'd2093733376, - 'd29720462, 'd65909788672, - 'd4543711744, - 'd2117079296, - 'd51891092, 'd67774132224, - 'd2911243008, - 'd2115622528, - 'd73113720, 'd68820041728, - 'd1273183616, - 'd2089790208, - 'd93158192, 'd69049499648, 'd351433280, - 'd2040284416, - 'd111811808, 'd68473896960, 'd1944049536, - 'd1968069376, - 'd128881496, 'd67113725952, 'd3486789120, - 'd1874356352, - 'd144195728, 'd64998219776, 'd4962652672, - 'd1760584960, - 'd157606112, 'd62164844544, 'd6355700736, - 'd1628403200, - 'd168988784, 'd58658750464, 'd7651218944, - 'd1479644416, - 'd178245392, 'd54532087808, 'd8835868672, - 'd1316303360, - 'd185303792, 'd49843318784, 'd9897820160, - 'd1140510208, - 'd190118496, 'd44656418816, 'd10826858496, - 'd954503680, - 'd192670752, 'd39040032768, 'd11614480384, - 'd760603392, - 'd192968256, 'd33066635264, 'd12253963264, - 'd561181504, - 'd191044672, 'd26811590656, 'd12740410368, - 'd358634592, - 'd186958800, 'd20352258048, 'd13070778368, - 'd155355344, - 'd180793488, 'd13767048192, 'd13243881472, 'd46295076, - 'd172654240, 'd7134508032, 'd13260374016, 'd244013680, - 'd162667648, 'd532402080, 'd13122712576, 'd435581472, - 'd150979568, - 'd5963171840, 'd12835095552, 'd618887680, - 'd137753088, - 'd12278635520, 'd12403388416, 'd791952384, - 'd123166384, - 'd18343737344, 'd11835023360, 'd952947136, - 'd107410400, - 'd24092315648, 'd11138892800, 'd1100213760, - 'd90686408, - 'd29462990848, 'd10325217280, 'd1232280576, - 'd73203528, - 'd34399793152, 'd9405405184, 'd1347876480, - 'd55176152, - 'd38852730880, 'd8391904768, 'd1445942016, - 'd36821416, - 'd42778251264, 'd7298036736, 'd1525638272, - 'd18356602, - 'd46139658240, 'd6137830912, 'd1586352896, 'd3364, - 'd48907403264, 'd4925849088, 'd1627703296, 'd18048354, - 'd51059314688, 'd3677007104, 'd1649537408, 'd35575396, - 'd52580737024, 'd2406398464, 'd1651931392, 'd52390896, - 'd53464559616, 'd1129114624, 'd1635185152, 'd68312728, - 'd53711183872, - 'd139928944, 'd1599814784, 'd83172152, - 'd53328396288, - 'd1386162304, 'd1546543488, 'd96815528, - 'd52331134976, - 'd2595524096, 'd1476289152, 'd109105848, - 'd50741219328, - 'd3754616064, 'd1390150784, 'd119924056, - 'd48586973184, - 'd4850846208, 'd1289392896, 'd129170104, - 'd45902774272, - 'd5872562688, 'd1175427840, 'd136763808, - 'd42728583168, - 'd6809170432, 'd1049796992, 'd142645424, - 'd39109353472, - 'd7651239424, 'd914150976, 'd146776032, - 'd35094458368, - 'd8390590464, 'd770228544, 'd149137584, - 'd30737025024, - 'd9020372992, 'd619834944, 'd149732832, - 'd26093264896, - 'd9535118336, 'd464820192, 'd148584864, - 'd21221765120, - 'd9930782720, 'd307056544, 'd145736576, - 'd16182777856, - 'd10204768256, 'd148416656, 'd141249808, - 'd11037487104, - 'd10355931136, - 'd9248055, 'd135204288, - 'd5847291392, - 'd10384567296, - 'd164128624, 'd127696448, - 'd673083584, - 'd10292387840, - 'd314478656, 'd118838032, 'd4425443328, - 'd10082473984, - 'd458633504, 'd108754496, 'd9390467072, - 'd9759219712, - 'd595028224, 'd97583376, 'd14166675456, - 'd9328256000, - 'd722214016, 'd85472480, 'd18701864960, - 'd8796367872, - 'd838872960, 'd72578000, 'd22947489792, - 'd8171397632, - 'd943831040, 'd59062548, 'd26859171840, - 'd7462130688, - 'd1036069504, 'd45093212, 'd30397132800, - 'd6678184448, - 'd1114734080, 'd30839494, 'd33526589440, - 'd5829879808, - 'd1179141760, 'd16471352, 'd36218060800, - 'd4928109056, - 'd1228786048, 'd2157196, 'd38447636480, - 'd3984203008, - 'd1263340160, - 'd11938022, 'd40197140480, - 'd3009790464, - 'd1282657280, - 'd25654662, 'd41454268416, - 'd2016659712, - 'd1286769408, - 'd38840152, 'd42212614144, - 'd1016618176, - 'd1275884288, - 'd51350640, 'd42471653376, - 'd21356334, - 'd1250379776, - 'd63052516, 'd42236645376, 'd957685888, - 'd1210796416, - 'd73823768, 'd41518489600, 'd1909447296, - 'd1157828864, - 'd83555224, 'd40333484032, 'd2823367424, - 'd1092315392, - 'd92151592, 'd38703067136, 'd3689500160, - 'd1015224960, - 'd99532312, 'd36653469696, 'd4498618368, - 'd927644736, - 'd105632264, 'd34215340032, 'd5242309120, - 'd830765056, - 'd110402272, 'd31423309824, 'd5913057792, - 'd725863872, - 'd113809368, 'd28315527168, 'd6504319488, - 'd614290688, - 'd115836928, 'd24933158912, 'd7010576896, - 'd497449664, - 'd116484592, 'd21319860224, 'd7427391488, - 'd376782464, - 'd115767992, 'd17521235968, 'd7751432704, - 'd253750912, - 'd113718288, 'd13584269312, 'd7980498432, - 'd129819680, - 'd110381560, 'd9556759552, 'd8113524224, - 'd6439408, - 'd105818040, 'd5486758400, 'd8150574080, 'd114969968, - 'd100101136, 'd1422006400, 'd8092821504, 'd233035072, - 'd93316416, - 'd2590614528, 'd7942518272, 'd346444256, - 'd85560352, - 'd6505608704, 'd7702948864, 'd453961664, - 'd76939064, - 'd10279368704, 'd7378376192, 'd554440448, - 'd67566928, - 'd13870651392, 'd6973975552, 'd646834304, - 'd57565096, - 'd17241012224, 'd6495759872, 'd730208128, - 'd47059976, - 'd20355205120, 'd5950494720, 'd803746816, - 'd36181704, - 'd23181537280, 'd5345609216, 'd866762944, - 'd25062552, - 'd25692176384, 'd4689098240, 'd918702144, - 'd13835381, - 'd27863408640, 'd3989420544, 'd959147840, - 'd2632072, - 'd29675841536, 'd3255392000, 'd987823232, 'd8417969, - 'd31114557440, 'd2496078848, 'd1004592512, 'd19189274, - 'd32169211904, 'd1720688896, 'd1009460096, 'd29561700, - 'd32834078720, 'd938460864, 'd1002568000, 'd39421732, - 'd33108035584, 'd158558640, 'd984192000, 'd48663680, - 'd32994498560, - 'd610034432, 'd954736192, 'd57190776};
endpackage
`endif
