`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam N = 2;
	localparam M = 2;
	localparam real Lfr[0:1] = {0.93051463, 0.93051463};
	localparam real Lfi[0:1] = {0.086347975, -0.086347975};
	localparam real Lbr[0:1] = {0.93051463, 0.93051463};
	localparam real Lbi[0:1] = {0.086347975, -0.086347975};
	localparam real Wfr[0:1] = {-0.011232297, -0.011232297};
	localparam real Wfi[0:1] = {-0.017049037, 0.017049037};
	localparam real Wbr[0:1] = {-0.011232297, -0.011232297};
	localparam real Wbi[0:1] = {-0.017049037, 0.017049037};
	localparam real Ffr[0:1][0:39] = '{
		'{-0.059192378, -0.24018086, -0.16673705, -0.20842467, -0.25860903, -0.17813122, -0.33566526, -0.14948735, -0.3988361, -0.12263594, -0.44910467, -0.09767976, -0.487488, -0.074685276, -0.5150203, -0.053686436, -0.53273803, -0.034688376, -0.54166687, -0.017670995, -0.5428106, -0.0025924132, -0.53714144, 0.0106077595, -0.5255922, 0.022005338, -0.5090496, 0.03168868, -0.4883494, 0.039756004, -0.4642727, 0.046312932, -0.437543, 0.051470272, -0.4088247, 0.055341974, -0.37872255, 0.058043353, -0.34778166, 0.059689485},
		'{-0.059192378, -0.24018086, -0.16673705, -0.20842467, -0.25860903, -0.17813122, -0.33566526, -0.14948735, -0.3988361, -0.12263594, -0.44910467, -0.09767976, -0.487488, -0.074685276, -0.5150203, -0.053686436, -0.53273803, -0.034688376, -0.54166687, -0.017670995, -0.5428106, -0.0025924132, -0.53714144, 0.0106077595, -0.5255922, 0.022005338, -0.5090496, 0.03168868, -0.4883494, 0.039756004, -0.4642727, 0.046312932, -0.437543, 0.051470272, -0.4088247, 0.055341974, -0.37872255, 0.058043353, -0.34778166, 0.059689485}};
	localparam real Ffi[0:1][0:39] = '{
		'{1.2931129, -0.1744933, 1.1981493, -0.1831077, 1.100498, -0.18838143, 1.0016991, -0.19067295, 0.90311164, -0.19033189, 0.8059199, -0.18769597, 0.71114093, -0.18308829, 0.61963344, -0.17681526, 0.532107, -0.1691649, 0.4491325, -0.16040568, 0.37115252, -0.15078568, 0.29849225, -0.14053212, 0.23137031, -0.12985124, 0.16990964, -0.11892836, 0.114148006, -0.10792832, 0.06404841, -0.09699603, 0.019508973, -0.0862572, -0.019627567, -0.075819224, -0.05356492, -0.06577223, -0.08254487, -0.056190096},
		'{-1.2931129, 0.1744933, -1.1981493, 0.1831077, -1.100498, 0.18838143, -1.0016991, 0.19067295, -0.90311164, 0.19033189, -0.8059199, 0.18769597, -0.71114093, 0.18308829, -0.61963344, 0.17681526, -0.532107, 0.1691649, -0.4491325, 0.16040568, -0.37115252, 0.15078568, -0.29849225, 0.14053212, -0.23137031, 0.12985124, -0.16990964, 0.11892836, -0.114148006, 0.10792832, -0.06404841, 0.09699603, -0.019508973, 0.0862572, 0.019627567, 0.075819224, 0.05356492, 0.06577223, 0.08254487, 0.056190096}};
	localparam real Fbr[0:1][0:39] = '{
		'{-0.059192378, 0.24018086, -0.16673705, 0.20842467, -0.25860903, 0.17813122, -0.33566526, 0.14948735, -0.3988361, 0.12263594, -0.44910467, 0.09767976, -0.487488, 0.074685276, -0.5150203, 0.053686436, -0.53273803, 0.034688376, -0.54166687, 0.017670995, -0.5428106, 0.0025924132, -0.53714144, -0.0106077595, -0.5255922, -0.022005338, -0.5090496, -0.03168868, -0.4883494, -0.039756004, -0.4642727, -0.046312932, -0.437543, -0.051470272, -0.4088247, -0.055341974, -0.37872255, -0.058043353, -0.34778166, -0.059689485},
		'{-0.059192378, 0.24018086, -0.16673705, 0.20842467, -0.25860903, 0.17813122, -0.33566526, 0.14948735, -0.3988361, 0.12263594, -0.44910467, 0.09767976, -0.487488, 0.074685276, -0.5150203, 0.053686436, -0.53273803, 0.034688376, -0.54166687, 0.017670995, -0.5428106, 0.0025924132, -0.53714144, -0.0106077595, -0.5255922, -0.022005338, -0.5090496, -0.03168868, -0.4883494, -0.039756004, -0.4642727, -0.046312932, -0.437543, -0.051470272, -0.4088247, -0.055341974, -0.37872255, -0.058043353, -0.34778166, -0.059689485}};
	localparam real Fbi[0:1][0:39] = '{
		'{1.2931129, 0.1744933, 1.1981493, 0.1831077, 1.100498, 0.18838143, 1.0016991, 0.19067295, 0.90311164, 0.19033189, 0.8059199, 0.18769597, 0.71114093, 0.18308829, 0.61963344, 0.17681526, 0.532107, 0.1691649, 0.4491325, 0.16040568, 0.37115252, 0.15078568, 0.29849225, 0.14053212, 0.23137031, 0.12985124, 0.16990964, 0.11892836, 0.114148006, 0.10792832, 0.06404841, 0.09699603, 0.019508973, 0.0862572, -0.019627567, 0.075819224, -0.05356492, 0.06577223, -0.08254487, 0.056190096},
		'{-1.2931129, -0.1744933, -1.1981493, -0.1831077, -1.100498, -0.18838143, -1.0016991, -0.19067295, -0.90311164, -0.19033189, -0.8059199, -0.18769597, -0.71114093, -0.18308829, -0.61963344, -0.17681526, -0.532107, -0.1691649, -0.4491325, -0.16040568, -0.37115252, -0.15078568, -0.29849225, -0.14053212, -0.23137031, -0.12985124, -0.16990964, -0.11892836, -0.114148006, -0.10792832, -0.06404841, -0.09699603, -0.019508973, -0.0862572, 0.019627567, -0.075819224, 0.05356492, -0.06577223, 0.08254487, -0.056190096}};
	localparam real hf[0:599] = {0.04542239, -0.0005543194, 0.04460026, -0.0015614439, 0.043334406, -0.0024217982, 0.041696593, -0.0031434074, 0.039754055, -0.003734984, 0.03756927, -0.0042057345, 0.035199758, -0.0045651835, 0.032698028, -0.004823015, 0.030111566, -0.0049889362, 0.027482878, -0.0050725527, 0.024849605, -0.0050832634, 0.022244675, -0.005030174, 0.019696496, -0.004922018, 0.017229183, -0.0047671013, 0.014862798, -0.00457325, 0.012613625, -0.004347779, 0.0104944445, -0.0040974626, 0.008514819, -0.0038285244, 0.0066813882, -0.0035466265, 0.004998153, -0.003256874, 0.0034667628, -0.0029638212, 0.0020867928, -0.002671486, 0.000856012, -0.0023833688, -0.00022936086, -0.0021024742, -0.001174414, -0.0018313382, -0.0019853148, -0.0015720549, -0.0026690974, -0.0013263079, -0.0032334663, -0.0010954011, -0.0036866167, -0.00088029105, -0.004037072, -0.00068161887, -0.004293537, -0.00049974263, -0.0044647683, -0.00033476876, -0.0045594615, -0.00018658249, -0.0045861485, -5.487742e-05, -0.004553118, 6.081651e-05, -0.0044683404, 0.0001611065, -0.004339413, 0.000246712, -0.0041735126, 0.0003184418, -0.0039773616, 0.0003771726, -0.0037572016, 0.0004238297, -0.0035187786, 0.0004593696, -0.0032673355, 0.00048476408, -0.00300761, 0.00050098647, -0.0027438423, 0.0005089995, -0.0024797847, 0.00050974474, -0.0022187172, 0.00050413376, -0.0019634685, 0.0004930408, -0.0017164368, 0.00047729647, -0.0014796156, 0.00045768355, -0.0012546206, 0.00043493308, -0.0010427174, 0.00040972198, -0.00084485055, 0.0003826717, -0.0006616725, 0.0003543475, -0.00049357256, 0.0003252587, -0.00034070548, 0.00029585956, -0.0002030193, 0.0002665505, -8.0282196e-05, 0.00023768011, 2.7891969e-05, 0.00020954752, 0.000122019286, 0.00018240484, 0.00020272304, 0.00015646007, 0.0002707124, 0.00013188018, 0.00032676294, 0.00010879418, 0.0003716986, 8.7296416e-05, 0.00040637553, 6.744977e-05, 0.00043166734, 4.928886e-05, 0.00044845234, 3.2823224e-05, 0.00045760203, 1.8040351e-05, 0.0004599713, 4.9086607e-06, 0.00045639006, -6.6197194e-06, 0.00044765612, -1.6606291e-05, 0.00043452956, -2.5123702e-05, 0.00041772812, -3.2253447e-05, 0.00039792372, -3.8083745e-05, 0.0003757401, -4.270759e-05, 0.00035175122, -4.622103e-05, 0.00032648043, -4.8721573e-05, 0.00030040054, -5.030683e-05, 0.00027393445, -5.1073275e-05, 0.0002474562, -5.111523e-05, 0.00022129256, -5.052396e-05, 0.00019572514, -4.9386945e-05, 0.00017099243, -4.77873e-05, 0.0001472925, -4.580328e-05, 0.00012478569, -4.3507953e-05, 0.00010359729, -4.0968953e-05, 8.382057e-05, -3.8248338e-05, 6.551963e-05, -3.540254e-05, 4.873231e-05, -3.2482374e-05, 3.3473083e-05, -2.9533136e-05, 1.973581e-05, -2.6594735e-05, 7.4964237e-06, -2.3701894e-05, -3.2844837e-06, -2.088438e-05, -1.2659248e-05, -1.8167259e-05, -2.0690846e-05, -1.5571191e-05, -2.7450777e-05, -1.311273e-05, -3.3017106e-05, -1.0804644e-05, -3.7472666e-05, -8.656235e-06, -4.0903447e-05, -6.673666e-06, -4.339713e-05, -4.8602815e-06, -4.5041794e-05, -3.2169237e-06, -4.59248e-05, -1.74224e-06, -4.613179e-05, -4.3297692e-07, -4.574587e-05, 7.157389e-07, -4.484689e-05, 1.7101355e-06, -4.3510885e-05, 2.5575478e-06, -4.1809642e-05, 3.266187e-06, -3.9810326e-05, 3.8449284e-06, -3.7575257e-05, 4.3031196e-06, -3.5161764e-05, 4.6504033e-06, -3.262209e-05, 4.896565e-06, -3.0003424e-05, 5.0513904e-06, -2.734794e-05, 5.1245493e-06, -2.4692923e-05, 5.125489e-06, -2.2070928e-05, 5.0633475e-06, -1.9509982e-05, 4.946879e-06, -1.7033808e-05, 4.7843973e-06, -1.4662086e-05, 4.5837273e-06, -1.2410717e-05, 4.3521723e-06, -1.0292111e-05, 4.096489e-06, -8.315474e-06, 3.8228754e-06, -6.4871015e-06, 3.5369642e-06, -4.81067e-06, 3.2438252e-06, -3.287525e-06, 2.9479752e-06, -1.9169574e-06, 2.653392e-06, -6.9647416e-07, 2.3635337e-06, 3.7794592e-07, 2.0813625e-06, 1.3116086e-06, 1.8093708e-06, 2.1108767e-06, 1.54961e-06, 2.7829578e-06, 1.3037219e-06, 3.335709e-06, 1.0729692e-06, 3.7774576e-06, 8.582693e-07, 4.116839e-06, 6.602258e-07, 4.3626537e-06, 4.7916143e-07, 4.5237357e-06, 3.1514938e-07, 4.60884e-06, 1.6804408e-07, 4.626547e-06, 3.7510784e-08, 4.5851766e-06, -7.6946485e-08, 4.492723e-06, -1.7595833e-07, 4.356792e-06, -2.602652e-07, 4.1845624e-06, -3.3069438e-07, 3.982748e-06, -3.881388e-07, 3.7575755e-06, -4.3353782e-07, 3.5147707e-06, -4.678597e-07, 3.25955e-06, -4.920862e-07, 2.9966213e-06, -5.0719865e-07, 2.7301912e-06, -5.1416606e-07, 2.463976e-06, -5.1393465e-07, 2.2012186e-06, -5.0741926e-07, 1.944709e-06, -4.9549607e-07, 1.6968066e-06, -4.7899664e-07, 1.4594661e-06, -4.5870337e-07, 1.2342651e-06, -4.3534615e-07, 1.0224321e-06, -4.0960015e-07, 8.248758e-07, -3.8208418e-07, 6.422143e-07, -3.5336055e-07, 4.7480444e-07, -3.2393504e-07, 3.2277057e-07, -2.942581e-07, 1.860324e-07, -2.6472605e-07, 6.433185e-08, -2.3568342e-07, -4.2741135e-08, -2.074249e-07, -1.3572436e-07, -1.8019833e-07, -2.1526061e-07, -1.5420738e-07, -2.8207637e-07, -1.2961485e-07, -3.369624e-07, -1.06545635e-07, -3.8075578e-07, -8.509016e-08, -4.1432386e-07, -6.530753e-08, -4.3854968e-07, -4.7228852e-08, -4.5431918e-07, -3.086033e-08, -4.6250995e-07, -1.618639e-08, -4.639815e-07, -3.1726002e-09, -4.59567e-07, 8.231488e-09, -4.5006632e-07, 1.8089715e-08, -4.3624058e-07, 2.6476819e-08, -4.188075e-07, 3.347614e-08, -3.9843823e-07, 3.9177518e-08, -3.75755e-07, 4.3675342e-08, -3.513296e-07, 4.7066838e-08, -3.2568275e-07, 4.9450495e-08, -2.9928427e-07, 5.092472e-08, -2.7255365e-07, 5.1586607e-08, -2.4586134e-07, 5.1530943e-08, -2.1953038e-07, 5.0849316e-08, -1.9383845e-07, 4.96294e-08, -1.6902018e-07, 4.7954373e-08, -1.452698e-07, 4.5902468e-08, -1.2274373e-07, 4.354664e-08, -1.01563614e-07, 4.0954323e-08, -8.181911e-08, 3.818733e-08, -6.357089e-08, 3.5301778e-08, -4.685355e-08, 3.2348133e-08, -3.1678518e-08, 2.9371304e-08, -1.8036815e-08, 2.6410795e-08, -5.9017635e-09, 2.350091e-08, 4.768437e-09, 2.0670978e-08, 1.40282905e-08, 1.7945634e-08, 2.1942718e-08, 1.5345107e-08, 2.8584946e-08, 1.2885529e-08, 3.403455e-08, 1.0579259e-08, 3.8375674e-08, 8.4352045e-09, 4.1695422e-08, 6.4591537e-09, 4.408241e-08, 4.654096e-09, 4.5625477e-08, 3.0205436e-09, 4.641259e-08, 1.5568352e-09, 4.6529845e-08, 2.5943456e-10, 4.6060663e-08, -8.7678975e-10, 4.5085102e-08, -1.8582991e-09, 4.3679297e-08, -2.6926366e-09, 4.1915026e-08, -3.388198e-09, 3.985937e-08, -3.95402e-09, 3.7574498e-08, -4.3995874e-09, 3.5117516e-08, -4.7346624e-09, 3.2540413e-08, -4.9691264e-09, 2.989006e-08, -5.1128453e-09, 2.7208294e-08, -5.1755493e-09, 2.4532042e-08, -5.166733e-09, 2.1893479e-08, -5.0955635e-09, 1.9320243e-08, -4.9708158e-09, 1.6835667e-08, -4.8008095e-09, 1.4459041e-08, -4.5933666e-09, 1.2205884e-08, -4.3557784e-09, 1.0088233e-08, -4.094782e-09, 8.114934e-09, -3.8165493e-09, 6.29194e-09, -3.5266816e-09, 4.622603e-09, -3.2302139e-09, 3.1079643e-09, -2.931624e-09, 1.747031e-09, -2.634849e-09, 5.370488e-10, -2.3433042e-09, -5.2624205e-10, -2.059909e-09, -1.4483639e-09, -1.7871115e-09, -2.235873e-09, -1.5269207e-09, -2.8961498e-09, -1.2809356e-09, -3.4372012e-09, -1.0503781e-09, -3.8674854e-09, -8.361263e-10, -4.1957495e-09, -6.387461e-10, -4.4308854e-09, -4.5852486e-10, -4.5818034e-09, -2.9550262e-10, -4.657318e-09, -1.4950312e-10, -4.6660547e-09, -2.0163262e-11, -4.6163655e-09, 9.303866e-11, -4.5162634e-09, 1.9075651e-10, -4.373364e-09, 2.7375152e-10, -4.1948445e-09, 3.4286937e-10, -3.9874113e-09, 3.9901904e-10, -3.7572745e-09, 4.4315368e-10, -3.5101382e-09, 4.7625326e-10, -3.2511915e-09, 4.993092e-10, -2.9851115e-09, 5.133106e-10, -2.7160707e-09, 5.1923266e-10, -2.447749e-09, 5.180261e-10, -2.1833513e-09, 5.106089e-10, -1.9256288e-09, 4.9785887e-10, -1.6769013e-09, 4.8060833e-10, -1.4390849e-09, 4.5963935e-10, -1.2137186e-09, 4.3568055e-10, -1.0019937e-09, 4.09405e-10, -8.047828e-10, 3.8142903e-10, -6.226698e-10, 3.5231165e-10, -4.5597906e-10, 3.2255523e-10, -3.0480446e-10, 2.926062e-10, -1.690374e-10, 2.6285688e-10, -4.8393695e-11, 2.336474e-10, 5.756054e-11, 2.0526823e-10, 1.4938471e-10, 1.7796276e-10, 2.2774092e-10, 1.5193038e-10, 2.9337283e-10, 1.2732963e-10, 3.4708622e-10, 1.0428132e-10, 3.8973116e-10, 8.2871904e-11, 4.2218604e-10, 6.3156765e-11, 4.453431e-10, 4.5163435e-11, 4.6009577e-10, 2.8894826e-11, 4.673276e-10, 1.433228e-11, 4.679025e-10, 1.4385536e-12, 4.6265677e-10, -9.839383e-12, 4.5239223e-10, -1.9567686e-11, 4.378708e-10, -2.782317e-11, 4.1981016e-10, -3.4691014e-11, 3.988805e-10, -4.026264e-11, 3.7570247e-10, -4.463382e-11, 3.5084555e-10, -4.7902942e-11, 3.2482783e-10, -5.0169462e-11, 2.9811595e-10, -5.1532553e-11, 2.71126e-10, -5.208992e-11, 2.4422475e-10, -5.1936795e-11, 2.1773142e-10, -5.116507e-11, 1.9191979e-10, -4.9862586e-11, 1.6702056e-10, -4.811259e-11, 1.4322403e-10, -4.599327e-11, 1.206828e-10, -4.357745e-11, 9.951475e-11, -4.093237e-11, 7.9805954e-11, -3.8119563e-11, 6.1613645e-11, -3.5194833e-11, 4.496918e-11, -3.2208288e-11, 2.9880938e-11, -2.9204444e-11, 1.6337112e-11, -2.6222394e-11, 4.3084178e-12, -2.329601e-11, -6.2493274e-12, -2.0454185e-11, -1.539278e-11, -1.772112e-11, -2.3188791e-11, -1.5116606e-11, -2.97123e-11, -1.2656355e-11, -3.5044374e-11, -1.0352312e-11};
	localparam real hb[0:599] = {0.04542239, 0.0005543194, 0.04460026, 0.0015614439, 0.043334406, 0.0024217982, 0.041696593, 0.0031434074, 0.039754055, 0.003734984, 0.03756927, 0.0042057345, 0.035199758, 0.0045651835, 0.032698028, 0.004823015, 0.030111566, 0.0049889362, 0.027482878, 0.0050725527, 0.024849605, 0.0050832634, 0.022244675, 0.005030174, 0.019696496, 0.004922018, 0.017229183, 0.0047671013, 0.014862798, 0.00457325, 0.012613625, 0.004347779, 0.0104944445, 0.0040974626, 0.008514819, 0.0038285244, 0.0066813882, 0.0035466265, 0.004998153, 0.003256874, 0.0034667628, 0.0029638212, 0.0020867928, 0.002671486, 0.000856012, 0.0023833688, -0.00022936086, 0.0021024742, -0.001174414, 0.0018313382, -0.0019853148, 0.0015720549, -0.0026690974, 0.0013263079, -0.0032334663, 0.0010954011, -0.0036866167, 0.00088029105, -0.004037072, 0.00068161887, -0.004293537, 0.00049974263, -0.0044647683, 0.00033476876, -0.0045594615, 0.00018658249, -0.0045861485, 5.487742e-05, -0.004553118, -6.081651e-05, -0.0044683404, -0.0001611065, -0.004339413, -0.000246712, -0.0041735126, -0.0003184418, -0.0039773616, -0.0003771726, -0.0037572016, -0.0004238297, -0.0035187786, -0.0004593696, -0.0032673355, -0.00048476408, -0.00300761, -0.00050098647, -0.0027438423, -0.0005089995, -0.0024797847, -0.00050974474, -0.0022187172, -0.00050413376, -0.0019634685, -0.0004930408, -0.0017164368, -0.00047729647, -0.0014796156, -0.00045768355, -0.0012546206, -0.00043493308, -0.0010427174, -0.00040972198, -0.00084485055, -0.0003826717, -0.0006616725, -0.0003543475, -0.00049357256, -0.0003252587, -0.00034070548, -0.00029585956, -0.0002030193, -0.0002665505, -8.0282196e-05, -0.00023768011, 2.7891969e-05, -0.00020954752, 0.000122019286, -0.00018240484, 0.00020272304, -0.00015646007, 0.0002707124, -0.00013188018, 0.00032676294, -0.00010879418, 0.0003716986, -8.7296416e-05, 0.00040637553, -6.744977e-05, 0.00043166734, -4.928886e-05, 0.00044845234, -3.2823224e-05, 0.00045760203, -1.8040351e-05, 0.0004599713, -4.9086607e-06, 0.00045639006, 6.6197194e-06, 0.00044765612, 1.6606291e-05, 0.00043452956, 2.5123702e-05, 0.00041772812, 3.2253447e-05, 0.00039792372, 3.8083745e-05, 0.0003757401, 4.270759e-05, 0.00035175122, 4.622103e-05, 0.00032648043, 4.8721573e-05, 0.00030040054, 5.030683e-05, 0.00027393445, 5.1073275e-05, 0.0002474562, 5.111523e-05, 0.00022129256, 5.052396e-05, 0.00019572514, 4.9386945e-05, 0.00017099243, 4.77873e-05, 0.0001472925, 4.580328e-05, 0.00012478569, 4.3507953e-05, 0.00010359729, 4.0968953e-05, 8.382057e-05, 3.8248338e-05, 6.551963e-05, 3.540254e-05, 4.873231e-05, 3.2482374e-05, 3.3473083e-05, 2.9533136e-05, 1.973581e-05, 2.6594735e-05, 7.4964237e-06, 2.3701894e-05, -3.2844837e-06, 2.088438e-05, -1.2659248e-05, 1.8167259e-05, -2.0690846e-05, 1.5571191e-05, -2.7450777e-05, 1.311273e-05, -3.3017106e-05, 1.0804644e-05, -3.7472666e-05, 8.656235e-06, -4.0903447e-05, 6.673666e-06, -4.339713e-05, 4.8602815e-06, -4.5041794e-05, 3.2169237e-06, -4.59248e-05, 1.74224e-06, -4.613179e-05, 4.3297692e-07, -4.574587e-05, -7.157389e-07, -4.484689e-05, -1.7101355e-06, -4.3510885e-05, -2.5575478e-06, -4.1809642e-05, -3.266187e-06, -3.9810326e-05, -3.8449284e-06, -3.7575257e-05, -4.3031196e-06, -3.5161764e-05, -4.6504033e-06, -3.262209e-05, -4.896565e-06, -3.0003424e-05, -5.0513904e-06, -2.734794e-05, -5.1245493e-06, -2.4692923e-05, -5.125489e-06, -2.2070928e-05, -5.0633475e-06, -1.9509982e-05, -4.946879e-06, -1.7033808e-05, -4.7843973e-06, -1.4662086e-05, -4.5837273e-06, -1.2410717e-05, -4.3521723e-06, -1.0292111e-05, -4.096489e-06, -8.315474e-06, -3.8228754e-06, -6.4871015e-06, -3.5369642e-06, -4.81067e-06, -3.2438252e-06, -3.287525e-06, -2.9479752e-06, -1.9169574e-06, -2.653392e-06, -6.9647416e-07, -2.3635337e-06, 3.7794592e-07, -2.0813625e-06, 1.3116086e-06, -1.8093708e-06, 2.1108767e-06, -1.54961e-06, 2.7829578e-06, -1.3037219e-06, 3.335709e-06, -1.0729692e-06, 3.7774576e-06, -8.582693e-07, 4.116839e-06, -6.602258e-07, 4.3626537e-06, -4.7916143e-07, 4.5237357e-06, -3.1514938e-07, 4.60884e-06, -1.6804408e-07, 4.626547e-06, -3.7510784e-08, 4.5851766e-06, 7.6946485e-08, 4.492723e-06, 1.7595833e-07, 4.356792e-06, 2.602652e-07, 4.1845624e-06, 3.3069438e-07, 3.982748e-06, 3.881388e-07, 3.7575755e-06, 4.3353782e-07, 3.5147707e-06, 4.678597e-07, 3.25955e-06, 4.920862e-07, 2.9966213e-06, 5.0719865e-07, 2.7301912e-06, 5.1416606e-07, 2.463976e-06, 5.1393465e-07, 2.2012186e-06, 5.0741926e-07, 1.944709e-06, 4.9549607e-07, 1.6968066e-06, 4.7899664e-07, 1.4594661e-06, 4.5870337e-07, 1.2342651e-06, 4.3534615e-07, 1.0224321e-06, 4.0960015e-07, 8.248758e-07, 3.8208418e-07, 6.422143e-07, 3.5336055e-07, 4.7480444e-07, 3.2393504e-07, 3.2277057e-07, 2.942581e-07, 1.860324e-07, 2.6472605e-07, 6.433185e-08, 2.3568342e-07, -4.2741135e-08, 2.074249e-07, -1.3572436e-07, 1.8019833e-07, -2.1526061e-07, 1.5420738e-07, -2.8207637e-07, 1.2961485e-07, -3.369624e-07, 1.06545635e-07, -3.8075578e-07, 8.509016e-08, -4.1432386e-07, 6.530753e-08, -4.3854968e-07, 4.7228852e-08, -4.5431918e-07, 3.086033e-08, -4.6250995e-07, 1.618639e-08, -4.639815e-07, 3.1726002e-09, -4.59567e-07, -8.231488e-09, -4.5006632e-07, -1.8089715e-08, -4.3624058e-07, -2.6476819e-08, -4.188075e-07, -3.347614e-08, -3.9843823e-07, -3.9177518e-08, -3.75755e-07, -4.3675342e-08, -3.513296e-07, -4.7066838e-08, -3.2568275e-07, -4.9450495e-08, -2.9928427e-07, -5.092472e-08, -2.7255365e-07, -5.1586607e-08, -2.4586134e-07, -5.1530943e-08, -2.1953038e-07, -5.0849316e-08, -1.9383845e-07, -4.96294e-08, -1.6902018e-07, -4.7954373e-08, -1.452698e-07, -4.5902468e-08, -1.2274373e-07, -4.354664e-08, -1.01563614e-07, -4.0954323e-08, -8.181911e-08, -3.818733e-08, -6.357089e-08, -3.5301778e-08, -4.685355e-08, -3.2348133e-08, -3.1678518e-08, -2.9371304e-08, -1.8036815e-08, -2.6410795e-08, -5.9017635e-09, -2.350091e-08, 4.768437e-09, -2.0670978e-08, 1.40282905e-08, -1.7945634e-08, 2.1942718e-08, -1.5345107e-08, 2.8584946e-08, -1.2885529e-08, 3.403455e-08, -1.0579259e-08, 3.8375674e-08, -8.4352045e-09, 4.1695422e-08, -6.4591537e-09, 4.408241e-08, -4.654096e-09, 4.5625477e-08, -3.0205436e-09, 4.641259e-08, -1.5568352e-09, 4.6529845e-08, -2.5943456e-10, 4.6060663e-08, 8.7678975e-10, 4.5085102e-08, 1.8582991e-09, 4.3679297e-08, 2.6926366e-09, 4.1915026e-08, 3.388198e-09, 3.985937e-08, 3.95402e-09, 3.7574498e-08, 4.3995874e-09, 3.5117516e-08, 4.7346624e-09, 3.2540413e-08, 4.9691264e-09, 2.989006e-08, 5.1128453e-09, 2.7208294e-08, 5.1755493e-09, 2.4532042e-08, 5.166733e-09, 2.1893479e-08, 5.0955635e-09, 1.9320243e-08, 4.9708158e-09, 1.6835667e-08, 4.8008095e-09, 1.4459041e-08, 4.5933666e-09, 1.2205884e-08, 4.3557784e-09, 1.0088233e-08, 4.094782e-09, 8.114934e-09, 3.8165493e-09, 6.29194e-09, 3.5266816e-09, 4.622603e-09, 3.2302139e-09, 3.1079643e-09, 2.931624e-09, 1.747031e-09, 2.634849e-09, 5.370488e-10, 2.3433042e-09, -5.2624205e-10, 2.059909e-09, -1.4483639e-09, 1.7871115e-09, -2.235873e-09, 1.5269207e-09, -2.8961498e-09, 1.2809356e-09, -3.4372012e-09, 1.0503781e-09, -3.8674854e-09, 8.361263e-10, -4.1957495e-09, 6.387461e-10, -4.4308854e-09, 4.5852486e-10, -4.5818034e-09, 2.9550262e-10, -4.657318e-09, 1.4950312e-10, -4.6660547e-09, 2.0163262e-11, -4.6163655e-09, -9.303866e-11, -4.5162634e-09, -1.9075651e-10, -4.373364e-09, -2.7375152e-10, -4.1948445e-09, -3.4286937e-10, -3.9874113e-09, -3.9901904e-10, -3.7572745e-09, -4.4315368e-10, -3.5101382e-09, -4.7625326e-10, -3.2511915e-09, -4.993092e-10, -2.9851115e-09, -5.133106e-10, -2.7160707e-09, -5.1923266e-10, -2.447749e-09, -5.180261e-10, -2.1833513e-09, -5.106089e-10, -1.9256288e-09, -4.9785887e-10, -1.6769013e-09, -4.8060833e-10, -1.4390849e-09, -4.5963935e-10, -1.2137186e-09, -4.3568055e-10, -1.0019937e-09, -4.09405e-10, -8.047828e-10, -3.8142903e-10, -6.226698e-10, -3.5231165e-10, -4.5597906e-10, -3.2255523e-10, -3.0480446e-10, -2.926062e-10, -1.690374e-10, -2.6285688e-10, -4.8393695e-11, -2.336474e-10, 5.756054e-11, -2.0526823e-10, 1.4938471e-10, -1.7796276e-10, 2.2774092e-10, -1.5193038e-10, 2.9337283e-10, -1.2732963e-10, 3.4708622e-10, -1.0428132e-10, 3.8973116e-10, -8.2871904e-11, 4.2218604e-10, -6.3156765e-11, 4.453431e-10, -4.5163435e-11, 4.6009577e-10, -2.8894826e-11, 4.673276e-10, -1.433228e-11, 4.679025e-10, -1.4385536e-12, 4.6265677e-10, 9.839383e-12, 4.5239223e-10, 1.9567686e-11, 4.378708e-10, 2.782317e-11, 4.1981016e-10, 3.4691014e-11, 3.988805e-10, 4.026264e-11, 3.7570247e-10, 4.463382e-11, 3.5084555e-10, 4.7902942e-11, 3.2482783e-10, 5.0169462e-11, 2.9811595e-10, 5.1532553e-11, 2.71126e-10, 5.208992e-11, 2.4422475e-10, 5.1936795e-11, 2.1773142e-10, 5.116507e-11, 1.9191979e-10, 4.9862586e-11, 1.6702056e-10, 4.811259e-11, 1.4322403e-10, 4.599327e-11, 1.206828e-10, 4.357745e-11, 9.951475e-11, 4.093237e-11, 7.9805954e-11, 3.8119563e-11, 6.1613645e-11, 3.5194833e-11, 4.496918e-11, 3.2208288e-11, 2.9880938e-11, 2.9204444e-11, 1.6337112e-11, 2.6222394e-11, 4.3084178e-12, 2.329601e-11, -6.2493274e-12, 2.0454185e-11, -1.539278e-11, 1.772112e-11, -2.3188791e-11, 1.5116606e-11, -2.97123e-11, 1.2656355e-11, -3.5044374e-11, 1.0352312e-11};
endpackage
`endif
