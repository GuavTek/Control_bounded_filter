`ifndef COEFFICIENTS_FX_SV_
`define COEFFICIENTS_FX_SV_

package Coefficients_Fx;

	localparam N = 4;
	localparam M = 4;
	localparam COEFF_BIAS = 48;
	localparam logic signed[63:0] Lfr[0:3] = {64'd275971144223279, 64'd275971144223279, 64'd270260315663771, 64'd270260315663771};

	localparam logic signed[63:0] Lfi[0:3] = {64'd22335262517471, - 64'd22335262517471, 64'd8848960108780, - 64'd8848960108780};

	localparam logic signed[63:0] Lbr[0:3] = {64'd275971144223279, 64'd275971144223279, 64'd270260315663771, 64'd270260315663771};

	localparam logic signed[63:0] Lbi[0:3] = {64'd22335262517471, - 64'd22335262517471, 64'd8848960108780, - 64'd8848960108780};

	localparam logic signed[63:0] Wfr[0:3] = {64'd28540176313, 64'd28540176313, 64'd8419923619, 64'd8419923619};

	localparam logic signed[63:0] Wfi[0:3] = {64'd1445518222, - 64'd1445518222, 64'd16512545571, - 64'd16512545571};

	localparam logic signed[63:0] Wbr[0:3] = {- 64'd28540176313, - 64'd28540176313, - 64'd8419923619, - 64'd8419923619};

	localparam logic signed[63:0] Wbi[0:3] = {- 64'd1445518222, 64'd1445518222, - 64'd16512545571, 64'd16512545571};

	localparam logic signed[63:0] Ffr[0:3][0:79] = '{
		'{64'd11318134054834866, 64'd1785088931865706, - 64'd339024165987731, 64'd6064496262143, 64'd12157123768699076, 64'd1570173789456536, - 64'd341272079255767, 64'd9172510400618, 64'd12887710479095196, 64'd1351740939832311, - 64'd341167778334080, 64'd12118475076591, 64'd13508529991771140, 64'd1131363344693918, - 64'd338788237891912, 64'd14887969489415, 64'd14018995473786920, 64'd910575946177082, - 64'd334223132521902, 64'd17468219104293, 64'd14419276164484444, 64'd690866648049596, - 64'd327573825977846, 64'd19848127586550, 64'd14710271727099088, 64'd473667903536096, - 64'd318952315119041, 64'd22018296491829, 64'd14893582553681816, 64'd260348946282488, - 64'd308480137083270, 64'd23971032977747, 64'd14971476352888860, 64'd52208695492740, - 64'd296287248179731, 64'd25700345873946, 64'd14946851364335296, - 64'd149530639238371, - 64'd282510882906723, 64'd27201930514309, 64'd14823196554594164, - 64'd343729233373810, - 64'd267294401359116, 64'd28473142797062, 64'd14604549158567508, - 64'd529334588597621, - 64'd250786133100118, 64'd29512962995340, 64'd14295449935890534, - 64'd705385730503098, - 64'd233138225333683, 64'd30321949892285, 64'd13900896515303776, - 64'd871016658879472, - 64'd214505502930986, 64'd30902185860766, 64'd13426295200604812, - 64'd1025459051789896, - 64'd195044347540348, 64'd31257213548188, 64'd12877411609950400, - 64'd1168044229578688, - 64'd174911602648054, 64'd31391964861468, 64'd12260320516016016, - 64'd1298204389689609, - 64'd154263511061512, 64'd31312682976210, 64'd11581355247939576, - 64'd1415473127694250, - 64'd133254690859766, 64'd31026838117143, 64'd10847057007198688, - 64'd1519485264197525, - 64'd112037155403479, 64'd30543037874340, 64'd10064124438726084, - 64'd1609976001285537, - 64'd90759382520839, 64'd29870932831370},
		'{64'd11318134054837492, 64'd1785088931865383, - 64'd339024165987741, 64'd6064496262145, 64'd12157123768701496, 64'd1570173789456241, - 64'd341272079255777, 64'd9172510400621, 64'd12887710479097400, 64'd1351740939832045, - 64'd341167778334089, 64'd12118475076593, 64'd13508529991773122, 64'd1131363344693683, - 64'd338788237891921, 64'd14887969489418, 64'd14018995473788672, 64'd910575946176876, - 64'd334223132521910, 64'd17468219104295, 64'd14419276164485964, 64'd690866648049422, - 64'd327573825977853, 64'd19848127586551, 64'd14710271727100368, 64'd473667903535953, - 64'd318952315119047, 64'd22018296491830, 64'd14893582553682860, 64'd260348946282376, - 64'd308480137083275, 64'd23971032977748, 64'd14971476352889670, 64'd52208695492659, - 64'd296287248179735, 64'd25700345873947, 64'd14946851364335868, - 64'd149530639238422, - 64'd282510882906727, 64'd27201930514310, 64'd14823196554594508, - 64'd343729233373832, - 64'd267294401359119, 64'd28473142797063, 64'd14604549158567628, - 64'd529334588597613, - 64'd250786133100121, 64'd29512962995341, 64'd14295449935890434, - 64'd705385730503062, - 64'd233138225333685, 64'd30321949892285, 64'd13900896515303468, - 64'd871016658879410, - 64'd214505502930987, 64'd30902185860766, 64'd13426295200604300, - 64'd1025459051789808, - 64'd195044347540347, 64'd31257213548187, 64'd12877411609949696, - 64'd1168044229578576, - 64'd174911602648054, 64'd31391964861468, 64'd12260320516015132, - 64'd1298204389689474, - 64'd154263511061511, 64'd31312682976209, 64'd11581355247938522, - 64'd1415473127694094, - 64'd133254690859764, 64'd31026838117142, 64'd10847057007197478, - 64'd1519485264197350, - 64'd112037155403476, 64'd30543037874339, 64'd10064124438724730, - 64'd1609976001285345, - 64'd90759382520835, 64'd29870932831369},
		'{64'd11105992628159936, 64'd1754361064338391, - 64'd315934402748876, 64'd73333543152989, 64'd11934023634477588, 64'd1559655744721768, - 64'd287263687069534, 64'd68836845288204, 64'd12667466654124698, 64'd1375946697860894, - 64'd260063825065816, 64'd64509577016534, 64'd13311726117986108, 64'd1202859200346066, - 64'd234291460699662, 64'd60349819761399, 64'd13872019441026244, 64'd1040020064829765, - 64'd209902904191354, 64'd56355371417979, 64'd14353378004129222, 64'd887058482823108, - 64'd186854270288440, 64'd52523773887942, 64'd14760648539409184, 64'd743606796377571, - 64'd165101606376356, 64'd48852339150369, 64'd15098494884311320, 64'd609301202147908, - 64'd144601010884036, 64'd45338173914597, 64'd15371400071548338, 64'd483782391236820, - 64'd125308742427901, 64'd41978202900829, 64'd15583668723593108, 64'd366696128125088, - 64'd107181320127219, 64'd38769190794348, 64'd15739429722075892, 64'd257693771893070, - 64'd90175615513249, 64'd35707762919080, 64'd15842639124012656, 64'd156432742840874, - 64'd74248936443612, 64'd32790424675987, 64'd15897083298320038, 64'd62576937515578, - 64'd59359103422214, 64'd30013579791484, 64'd15906382257551964, - 64'd24202904945215, - 64'd45464518713761, 64'd27373547420614, 64'd15873993161222760, - 64'd104228882343164, - 64'd32524228630416, 64'd24866578149255, 64'd15803213968462104, - 64'd177815652110490, - 64'd20497979356684, 64'd22488868939019, 64'd15697187219078688, - 64'd245270194548944, - 64'd9346266666974, 64'd20236577057897, 64'd15558903923391864, - 64'd306891614099658, 64'd969620121281, 64'd18105833038948, 64'd15391207542425108, - 64'd362970976223260, 64'd10487559627672, 64'd16092752708634, 64'd15196798041241474, - 64'd413791177564508, 64'd19244565002294, 64'd14193448325528},
		'{64'd11105992628167634, 64'd1754361064337296, - 64'd315934402748889, 64'd73333543152995, 64'd11934023634484916, 64'd1559655744720725, - 64'd287263687069546, 64'd68836845288210, 64'd12667466654131670, 64'd1375946697859902, - 64'd260063825065827, 64'd64509577016539, 64'd13311726117992736, 64'd1202859200345124, - 64'd234291460699673, 64'd60349819761404, 64'd13872019441032534, 64'd1040020064828870, - 64'd209902904191364, 64'd56355371417984, 64'd14353378004135182, 64'd887058482822260, - 64'd186854270288450, 64'd52523773887947, 64'd14760648539414826, 64'd743606796376768, - 64'd165101606376365, 64'd48852339150374, 64'd15098494884316656, 64'd609301202147149, - 64'd144601010884045, 64'd45338173914602, 64'd15371400071553376, 64'd483782391236103, - 64'd125308742427910, 64'd41978202900833, 64'd15583668723597856, 64'd366696128124412, - 64'd107181320127227, 64'd38769190794352, 64'd15739429722080360, 64'd257693771892434, - 64'd90175615513257, 64'd35707762919083, 64'd15842639124016860, 64'd156432742840275, - 64'd74248936443618, 64'd32790424675990, 64'd15897083298323982, 64'd62576937515016, - 64'd59359103422221, 64'd30013579791487, 64'd15906382257555660, - 64'd24202904945742, - 64'd45464518713767, 64'd27373547420617, 64'd15873993161226216, - 64'd104228882343657, - 64'd32524228630422, 64'd24866578149258, 64'd15803213968465330, - 64'd177815652110950, - 64'd20497979356689, 64'd22488868939022, 64'd15697187219081696, - 64'd245270194549373, - 64'd9346266666979, 64'd20236577057899, 64'd15558903923394660, - 64'd306891614100056, 64'd969620121277, 64'd18105833038950, 64'd15391207542427704, - 64'd362970976223631, 64'd10487559627668, 64'd16092752708636, 64'd15196798041243876, - 64'd413791177564851, 64'd19244565002290, 64'd14193448325529}};

	localparam logic signed[63:0] Ffi[0:3][0:79] = '{
		'{- 64'd13362176685608098, 64'd2268538559092143, 64'd111870794067565, - 64'd40662435826780, - 64'd12202795907676822, 64'd2365828819170948, 64'd82781487609260, - 64'd39386118636639, - 64'd10999510630446128, 64'd2444163023257960, 64'd54082606396732, - 64'd37888134581454, - 64'd9761781206594062, 64'd2503632696514646, 64'd25953166294419, - 64'd36185676786653, - 64'd8498991255300306, 64'd2544452390219278, - 64'd1437425228302, - 64'd34296746493141, - 64'd7220387478421469, 64'd2566954259288082, - 64'd27930188967951, - 64'd32240006623286, - 64'd5935022342774702, 64'd2571582030175910, - 64'd53377297621628, - 64'd30034635676189, - 64'd4651699918405561, 64'd2558884419213031, - 64'd77642701473218, - 64'd27700182917395, - 64'd3378925132237505, 64'd2529508063157622, - 64'd100602655128522, - 64'd25256425788224, - 64'd2124856665277585, 64'd2484190024997960, - 64'd122146144990124, - 64'd22723230415103, - 64'd897263689818794, 64'd2423749938831142, - 64'd142175217835754, - 64'd20120416050013, 64'd296513388937731, 64'd2349081857985880, - 64'd160605211512651, - 64'd17467624219949, 64'd1449598054494282, 64'd2261145870458153, - 64'd177364889381340, - 64'd14784193306640, 64'd2555608563476537, 64'd2160959545204884, - 64'd192396480732131, - 64'd12089039218089, 64'd3608684523992682, 64'd2049589271909884, - 64'd205655629953527, - 64'd9400542751380, 64'd4603509130055544, 64'd1928141555517314, - 64'd217111257751045, - 64'd6736444182049, 64'd5535327044432556, 64'd1797754325142296, - 64'd226745338195426, - 64'd4113745549702, 64'd6399957951599597, 64'd1659588314939304, - 64'd234552595818768, - 64'd1548621042939, 64'd7193805830690683, 64'd1514818572161070, - 64'd240540127374385, 64'd943664180559, 64'd7913864025303378, 64'd1364626145000200, - 64'd244726953229594, 64'd3348826470087},
		'{64'd13362176685606148, - 64'd2268538559091868, - 64'd111870794067560, 64'd40662435826778, 64'd12202795907674702, - 64'd2365828819170652, - 64'd82781487609254, 64'd39386118636637, 64'd10999510630443858, - 64'd2444163023257646, - 64'd54082606396726, 64'd37888134581452, 64'd9761781206591662, - 64'd2503632696514318, - 64'd25953166294412, 64'd36185676786650, 64'd8498991255297795, - 64'd2544452390218938, 64'd1437425228309, 64'd34296746493138, 64'd7220387478418869, - 64'd2566954259287732, 64'd27930188967959, 64'd32240006623283, 64'd5935022342772032, - 64'd2571582030175553, 64'd53377297621637, 64'd30034635676186, 64'd4651699918402839, - 64'd2558884419212670, 64'd77642701473226, 64'd27700182917392, 64'd3378925132234753, - 64'd2529508063157258, 64'd100602655128530, 64'd25256425788221, 64'd2124856665274824, - 64'd2484190024997598, 64'd122146144990133, 64'd22723230415101, 64'd897263689816041, - 64'd2423749938830783, 64'd142175217835764, 64'd20120416050010, - 64'd296513388940456, - 64'd2349081857985526, 64'd160605211512660, 64'd17467624219947, - 64'd1449598054496964, - 64'd2261145870457806, 64'd177364889381349, 64'd14784193306637, - 64'd2555608563479158, - 64'd2160959545204546, 64'd192396480732141, 64'd12089039218086, - 64'd3608684523995228, - 64'd2049589271909558, 64'd205655629953536, 64'd9400542751377, - 64'd4603509130057998, - 64'd1928141555517001, 64'd217111257751054, 64'd6736444182046, - 64'd5535327044434908, - 64'd1797754325141999, 64'd226745338195434, 64'd4113745549700, - 64'd6399957951601832, - 64'd1659588314939024, 64'd234552595818777, 64'd1548621042936, - 64'd7193805830692790, - 64'd1514818572160807, 64'd240540127374393, - 64'd943664180561, - 64'd7913864025305348, - 64'd1364626144999956, 64'd244726953229602, - 64'd3348826470089},
		'{- 64'd40413782719866184, 64'd3969970503004833, - 64'd511584607975589, 64'd50095953816924, - 64'd38454449186897512, 64'd3866950324012459, - 64'd501134098013000, 64'd50405453642227, - 64'd36547148869376472, 64'd3761913613303843, - 64'd490198617436206, 64'd50561255841662, - 64'd34692782275225136, 64'd3655286413364360, - 64'd478843729112543, 64'd50574810607094, - 64'd32892044130362836, 64'd3547466011602596, - 64'd467131020702752, 64'd50457051610484, - 64'd31145437456944600, 64'd3438822134314362, - 64'd455118252550944, 64'd50218407669809, - 64'd29453287059820696, 64'd3329698119571906, - 64'd442859504029156, 64'd49868814815822, - 64'd27815752432111084, 64'd3220412067642288, - 64'd430405318078685, 64'd49417728697649, - 64'd26232840091444668, 64'd3111257967704472, - 64'd417802843714956, 64'd48874137269154, - 64'd24704415358989096, 64'd3002506799790498, - 64'd405095976285888, 64'd48246573701731, - 64'd23230213593897208, 64'd2894407611022914, - 64'd392325495295720, 64'd47543129472821, - 64'd21809850896225256, 64'd2787188565358304, - 64'd379529199627015, 64'd46771467582875, - 64'd20442834291740392, 64'd2681057966175946, - 64'd366742040013165, 64'd45938835856821, - 64'd19128571412335052, 64'd2576205251171553, - 64'd353996248632204, 64'd45052080289263, - 64'd17866379686007044, 64'd2472801959129038, - 64'd341321465710084, 64'd44117658395658, - 64'd16655495050551182, 64'd2371002668248560, - 64'd328744863037924, 64'd43141652534621, - 64'd15495080205244352, 64'd2270945905807252, - 64'd316291264323036, 64'd42129783169274, - 64'd14384232414894556, 64'd2172755029020048, - 64'd303983262307876, 64'd41087422038180, - 64'd13321990880669480, 64'd2076539077052488, - 64'd291841332604490, 64'd40019605208908, - 64'd12307343692124342, 64'd1982393594215338, - 64'd279883944204475, 64'd38931045989650},
		'{64'd40413782719864280, - 64'd3969970503004567, 64'd511584607975594, - 64'd50095953816926, 64'd38454449186895440, - 64'd3866950324012170, 64'd501134098013006, - 64'd50405453642228, 64'd36547148869374256, - 64'd3761913613303532, 64'd490198617436211, - 64'd50561255841664, 64'd34692782275222784, - 64'd3655286413364030, 64'd478843729112549, - 64'd50574810607096, 64'd32892044130360372, - 64'd3547466011602249, 64'd467131020702757, - 64'd50457051610486, 64'd31145437456942032, - 64'd3438822134314002, 64'd455118252550949, - 64'd50218407669811, 64'd29453287059818048, - 64'd3329698119571532, 64'd442859504029161, - 64'd49868814815824, 64'd27815752432108364, - 64'd3220412067641905, 64'd430405318078690, - 64'd49417728697652, 64'd26232840091441888, - 64'd3111257967704080, 64'd417802843714961, - 64'd48874137269156, 64'd24704415358986264, - 64'd3002506799790098, 64'd405095976285894, - 64'd48246573701733, 64'd23230213593894340, - 64'd2894407611022510, 64'd392325495295726, - 64'd47543129472823, 64'd21809850896222364, - 64'd2787188565357896, 64'd379529199627020, - 64'd46771467582877, 64'd20442834291737480, - 64'd2681057966175535, 64'd366742040013170, - 64'd45938835856823, 64'd19128571412332136, - 64'd2576205251171141, 64'd353996248632210, - 64'd45052080289266, 64'd17866379686004130, - 64'd2472801959128626, 64'd341321465710090, - 64'd44117658395661, 64'd16655495050548274, - 64'd2371002668248148, 64'd328744863037930, - 64'd43141652534624, 64'd15495080205241458, - 64'd2270945905806842, 64'd316291264323041, - 64'd42129783169276, 64'd14384232414891682, - 64'd2172755029019642, 64'd303983262307882, - 64'd41087422038183, 64'd13321990880666632, - 64'd2076539077052086, 64'd291841332604495, - 64'd40019605208911, 64'd12307343692121528, - 64'd1982393594214940, 64'd279883944204480, - 64'd38931045989652}};

	localparam logic signed[63:0] Fbr[0:3][0:79] = '{
		'{- 64'd11318134054834866, 64'd1785088931865706, 64'd339024165987731, 64'd6064496262143, - 64'd12157123768699076, 64'd1570173789456536, 64'd341272079255767, 64'd9172510400618, - 64'd12887710479095196, 64'd1351740939832311, 64'd341167778334080, 64'd12118475076591, - 64'd13508529991771140, 64'd1131363344693918, 64'd338788237891912, 64'd14887969489415, - 64'd14018995473786920, 64'd910575946177082, 64'd334223132521902, 64'd17468219104293, - 64'd14419276164484444, 64'd690866648049596, 64'd327573825977846, 64'd19848127586550, - 64'd14710271727099088, 64'd473667903536096, 64'd318952315119041, 64'd22018296491829, - 64'd14893582553681816, 64'd260348946282488, 64'd308480137083270, 64'd23971032977747, - 64'd14971476352888860, 64'd52208695492740, 64'd296287248179731, 64'd25700345873946, - 64'd14946851364335296, - 64'd149530639238371, 64'd282510882906723, 64'd27201930514309, - 64'd14823196554594164, - 64'd343729233373810, 64'd267294401359116, 64'd28473142797062, - 64'd14604549158567508, - 64'd529334588597621, 64'd250786133100118, 64'd29512962995340, - 64'd14295449935890534, - 64'd705385730503098, 64'd233138225333683, 64'd30321949892285, - 64'd13900896515303776, - 64'd871016658879472, 64'd214505502930986, 64'd30902185860766, - 64'd13426295200604812, - 64'd1025459051789896, 64'd195044347540348, 64'd31257213548188, - 64'd12877411609950400, - 64'd1168044229578688, 64'd174911602648054, 64'd31391964861468, - 64'd12260320516016016, - 64'd1298204389689609, 64'd154263511061512, 64'd31312682976210, - 64'd11581355247939576, - 64'd1415473127694250, 64'd133254690859766, 64'd31026838117143, - 64'd10847057007198688, - 64'd1519485264197525, 64'd112037155403479, 64'd30543037874340, - 64'd10064124438726084, - 64'd1609976001285537, 64'd90759382520839, 64'd29870932831370},
		'{- 64'd11318134054837492, 64'd1785088931865383, 64'd339024165987741, 64'd6064496262145, - 64'd12157123768701496, 64'd1570173789456241, 64'd341272079255777, 64'd9172510400621, - 64'd12887710479097400, 64'd1351740939832045, 64'd341167778334089, 64'd12118475076593, - 64'd13508529991773122, 64'd1131363344693683, 64'd338788237891921, 64'd14887969489418, - 64'd14018995473788672, 64'd910575946176876, 64'd334223132521910, 64'd17468219104295, - 64'd14419276164485964, 64'd690866648049422, 64'd327573825977853, 64'd19848127586551, - 64'd14710271727100368, 64'd473667903535953, 64'd318952315119047, 64'd22018296491830, - 64'd14893582553682860, 64'd260348946282376, 64'd308480137083275, 64'd23971032977748, - 64'd14971476352889670, 64'd52208695492659, 64'd296287248179735, 64'd25700345873947, - 64'd14946851364335868, - 64'd149530639238422, 64'd282510882906727, 64'd27201930514310, - 64'd14823196554594508, - 64'd343729233373832, 64'd267294401359119, 64'd28473142797063, - 64'd14604549158567628, - 64'd529334588597613, 64'd250786133100121, 64'd29512962995341, - 64'd14295449935890434, - 64'd705385730503062, 64'd233138225333685, 64'd30321949892285, - 64'd13900896515303468, - 64'd871016658879410, 64'd214505502930987, 64'd30902185860766, - 64'd13426295200604300, - 64'd1025459051789808, 64'd195044347540347, 64'd31257213548187, - 64'd12877411609949696, - 64'd1168044229578576, 64'd174911602648054, 64'd31391964861468, - 64'd12260320516015132, - 64'd1298204389689474, 64'd154263511061511, 64'd31312682976209, - 64'd11581355247938522, - 64'd1415473127694094, 64'd133254690859764, 64'd31026838117142, - 64'd10847057007197478, - 64'd1519485264197350, 64'd112037155403476, 64'd30543037874339, - 64'd10064124438724730, - 64'd1609976001285345, 64'd90759382520835, 64'd29870932831369},
		'{- 64'd11105992628159936, 64'd1754361064338391, 64'd315934402748876, 64'd73333543152989, - 64'd11934023634477588, 64'd1559655744721768, 64'd287263687069534, 64'd68836845288204, - 64'd12667466654124698, 64'd1375946697860894, 64'd260063825065816, 64'd64509577016534, - 64'd13311726117986108, 64'd1202859200346066, 64'd234291460699662, 64'd60349819761399, - 64'd13872019441026244, 64'd1040020064829765, 64'd209902904191354, 64'd56355371417979, - 64'd14353378004129222, 64'd887058482823108, 64'd186854270288440, 64'd52523773887942, - 64'd14760648539409184, 64'd743606796377571, 64'd165101606376356, 64'd48852339150369, - 64'd15098494884311320, 64'd609301202147908, 64'd144601010884036, 64'd45338173914597, - 64'd15371400071548338, 64'd483782391236820, 64'd125308742427901, 64'd41978202900829, - 64'd15583668723593108, 64'd366696128125088, 64'd107181320127219, 64'd38769190794348, - 64'd15739429722075892, 64'd257693771893070, 64'd90175615513249, 64'd35707762919080, - 64'd15842639124012656, 64'd156432742840874, 64'd74248936443612, 64'd32790424675987, - 64'd15897083298320038, 64'd62576937515578, 64'd59359103422214, 64'd30013579791484, - 64'd15906382257551964, - 64'd24202904945215, 64'd45464518713761, 64'd27373547420614, - 64'd15873993161222760, - 64'd104228882343164, 64'd32524228630416, 64'd24866578149255, - 64'd15803213968462104, - 64'd177815652110490, 64'd20497979356684, 64'd22488868939019, - 64'd15697187219078688, - 64'd245270194548944, 64'd9346266666974, 64'd20236577057897, - 64'd15558903923391864, - 64'd306891614099658, - 64'd969620121281, 64'd18105833038948, - 64'd15391207542425108, - 64'd362970976223260, - 64'd10487559627672, 64'd16092752708634, - 64'd15196798041241474, - 64'd413791177564508, - 64'd19244565002294, 64'd14193448325528},
		'{- 64'd11105992628167634, 64'd1754361064337296, 64'd315934402748889, 64'd73333543152995, - 64'd11934023634484916, 64'd1559655744720725, 64'd287263687069546, 64'd68836845288210, - 64'd12667466654131670, 64'd1375946697859902, 64'd260063825065827, 64'd64509577016539, - 64'd13311726117992736, 64'd1202859200345124, 64'd234291460699673, 64'd60349819761404, - 64'd13872019441032534, 64'd1040020064828870, 64'd209902904191364, 64'd56355371417984, - 64'd14353378004135182, 64'd887058482822260, 64'd186854270288450, 64'd52523773887947, - 64'd14760648539414826, 64'd743606796376768, 64'd165101606376365, 64'd48852339150374, - 64'd15098494884316656, 64'd609301202147149, 64'd144601010884045, 64'd45338173914602, - 64'd15371400071553376, 64'd483782391236103, 64'd125308742427910, 64'd41978202900833, - 64'd15583668723597856, 64'd366696128124412, 64'd107181320127227, 64'd38769190794352, - 64'd15739429722080360, 64'd257693771892434, 64'd90175615513257, 64'd35707762919083, - 64'd15842639124016860, 64'd156432742840275, 64'd74248936443618, 64'd32790424675990, - 64'd15897083298323982, 64'd62576937515016, 64'd59359103422221, 64'd30013579791487, - 64'd15906382257555660, - 64'd24202904945742, 64'd45464518713767, 64'd27373547420617, - 64'd15873993161226216, - 64'd104228882343657, 64'd32524228630422, 64'd24866578149258, - 64'd15803213968465330, - 64'd177815652110950, 64'd20497979356689, 64'd22488868939022, - 64'd15697187219081696, - 64'd245270194549373, 64'd9346266666979, 64'd20236577057899, - 64'd15558903923394660, - 64'd306891614100056, - 64'd969620121277, 64'd18105833038950, - 64'd15391207542427704, - 64'd362970976223631, - 64'd10487559627668, 64'd16092752708636, - 64'd15196798041243876, - 64'd413791177564851, - 64'd19244565002290, 64'd14193448325529}};

	localparam logic signed[63:0] Fbi[0:3][0:79] = '{
		'{64'd13362176685608098, 64'd2268538559092143, - 64'd111870794067565, - 64'd40662435826780, 64'd12202795907676822, 64'd2365828819170948, - 64'd82781487609260, - 64'd39386118636639, 64'd10999510630446128, 64'd2444163023257960, - 64'd54082606396732, - 64'd37888134581454, 64'd9761781206594062, 64'd2503632696514646, - 64'd25953166294419, - 64'd36185676786653, 64'd8498991255300306, 64'd2544452390219278, 64'd1437425228302, - 64'd34296746493141, 64'd7220387478421469, 64'd2566954259288082, 64'd27930188967951, - 64'd32240006623286, 64'd5935022342774702, 64'd2571582030175910, 64'd53377297621628, - 64'd30034635676189, 64'd4651699918405561, 64'd2558884419213031, 64'd77642701473218, - 64'd27700182917395, 64'd3378925132237505, 64'd2529508063157622, 64'd100602655128522, - 64'd25256425788224, 64'd2124856665277585, 64'd2484190024997960, 64'd122146144990124, - 64'd22723230415103, 64'd897263689818794, 64'd2423749938831142, 64'd142175217835754, - 64'd20120416050013, - 64'd296513388937731, 64'd2349081857985880, 64'd160605211512651, - 64'd17467624219949, - 64'd1449598054494282, 64'd2261145870458153, 64'd177364889381340, - 64'd14784193306640, - 64'd2555608563476537, 64'd2160959545204884, 64'd192396480732131, - 64'd12089039218089, - 64'd3608684523992682, 64'd2049589271909884, 64'd205655629953527, - 64'd9400542751380, - 64'd4603509130055544, 64'd1928141555517314, 64'd217111257751045, - 64'd6736444182049, - 64'd5535327044432556, 64'd1797754325142296, 64'd226745338195426, - 64'd4113745549702, - 64'd6399957951599597, 64'd1659588314939304, 64'd234552595818768, - 64'd1548621042939, - 64'd7193805830690683, 64'd1514818572161070, 64'd240540127374385, 64'd943664180559, - 64'd7913864025303378, 64'd1364626145000200, 64'd244726953229594, 64'd3348826470087},
		'{- 64'd13362176685606148, - 64'd2268538559091868, 64'd111870794067560, 64'd40662435826778, - 64'd12202795907674702, - 64'd2365828819170652, 64'd82781487609254, 64'd39386118636637, - 64'd10999510630443858, - 64'd2444163023257646, 64'd54082606396726, 64'd37888134581452, - 64'd9761781206591662, - 64'd2503632696514318, 64'd25953166294412, 64'd36185676786650, - 64'd8498991255297795, - 64'd2544452390218938, - 64'd1437425228309, 64'd34296746493138, - 64'd7220387478418869, - 64'd2566954259287732, - 64'd27930188967959, 64'd32240006623283, - 64'd5935022342772032, - 64'd2571582030175553, - 64'd53377297621637, 64'd30034635676186, - 64'd4651699918402839, - 64'd2558884419212670, - 64'd77642701473226, 64'd27700182917392, - 64'd3378925132234753, - 64'd2529508063157258, - 64'd100602655128530, 64'd25256425788221, - 64'd2124856665274824, - 64'd2484190024997598, - 64'd122146144990133, 64'd22723230415101, - 64'd897263689816041, - 64'd2423749938830783, - 64'd142175217835764, 64'd20120416050010, 64'd296513388940456, - 64'd2349081857985526, - 64'd160605211512660, 64'd17467624219947, 64'd1449598054496964, - 64'd2261145870457806, - 64'd177364889381349, 64'd14784193306637, 64'd2555608563479158, - 64'd2160959545204546, - 64'd192396480732141, 64'd12089039218086, 64'd3608684523995228, - 64'd2049589271909558, - 64'd205655629953536, 64'd9400542751377, 64'd4603509130057998, - 64'd1928141555517001, - 64'd217111257751054, 64'd6736444182046, 64'd5535327044434908, - 64'd1797754325141999, - 64'd226745338195434, 64'd4113745549700, 64'd6399957951601832, - 64'd1659588314939024, - 64'd234552595818777, 64'd1548621042936, 64'd7193805830692790, - 64'd1514818572160807, - 64'd240540127374393, - 64'd943664180561, 64'd7913864025305348, - 64'd1364626144999956, - 64'd244726953229602, - 64'd3348826470089},
		'{64'd40413782719866184, 64'd3969970503004833, 64'd511584607975589, 64'd50095953816924, 64'd38454449186897512, 64'd3866950324012459, 64'd501134098013000, 64'd50405453642227, 64'd36547148869376472, 64'd3761913613303843, 64'd490198617436206, 64'd50561255841662, 64'd34692782275225136, 64'd3655286413364360, 64'd478843729112543, 64'd50574810607094, 64'd32892044130362836, 64'd3547466011602596, 64'd467131020702752, 64'd50457051610484, 64'd31145437456944600, 64'd3438822134314362, 64'd455118252550944, 64'd50218407669809, 64'd29453287059820696, 64'd3329698119571906, 64'd442859504029156, 64'd49868814815822, 64'd27815752432111084, 64'd3220412067642288, 64'd430405318078685, 64'd49417728697649, 64'd26232840091444668, 64'd3111257967704472, 64'd417802843714956, 64'd48874137269154, 64'd24704415358989096, 64'd3002506799790498, 64'd405095976285888, 64'd48246573701731, 64'd23230213593897208, 64'd2894407611022914, 64'd392325495295720, 64'd47543129472821, 64'd21809850896225256, 64'd2787188565358304, 64'd379529199627015, 64'd46771467582875, 64'd20442834291740392, 64'd2681057966175946, 64'd366742040013165, 64'd45938835856821, 64'd19128571412335052, 64'd2576205251171553, 64'd353996248632204, 64'd45052080289263, 64'd17866379686007044, 64'd2472801959129038, 64'd341321465710084, 64'd44117658395658, 64'd16655495050551182, 64'd2371002668248560, 64'd328744863037924, 64'd43141652534621, 64'd15495080205244352, 64'd2270945905807252, 64'd316291264323036, 64'd42129783169274, 64'd14384232414894556, 64'd2172755029020048, 64'd303983262307876, 64'd41087422038180, 64'd13321990880669480, 64'd2076539077052488, 64'd291841332604490, 64'd40019605208908, 64'd12307343692124342, 64'd1982393594215338, 64'd279883944204475, 64'd38931045989650},
		'{- 64'd40413782719864280, - 64'd3969970503004567, - 64'd511584607975594, - 64'd50095953816926, - 64'd38454449186895440, - 64'd3866950324012170, - 64'd501134098013006, - 64'd50405453642228, - 64'd36547148869374256, - 64'd3761913613303532, - 64'd490198617436211, - 64'd50561255841664, - 64'd34692782275222784, - 64'd3655286413364030, - 64'd478843729112549, - 64'd50574810607096, - 64'd32892044130360372, - 64'd3547466011602249, - 64'd467131020702757, - 64'd50457051610486, - 64'd31145437456942032, - 64'd3438822134314002, - 64'd455118252550949, - 64'd50218407669811, - 64'd29453287059818048, - 64'd3329698119571532, - 64'd442859504029161, - 64'd49868814815824, - 64'd27815752432108364, - 64'd3220412067641905, - 64'd430405318078690, - 64'd49417728697652, - 64'd26232840091441888, - 64'd3111257967704080, - 64'd417802843714961, - 64'd48874137269156, - 64'd24704415358986264, - 64'd3002506799790098, - 64'd405095976285894, - 64'd48246573701733, - 64'd23230213593894340, - 64'd2894407611022510, - 64'd392325495295726, - 64'd47543129472823, - 64'd21809850896222364, - 64'd2787188565357896, - 64'd379529199627020, - 64'd46771467582877, - 64'd20442834291737480, - 64'd2681057966175535, - 64'd366742040013170, - 64'd45938835856823, - 64'd19128571412332136, - 64'd2576205251171141, - 64'd353996248632210, - 64'd45052080289266, - 64'd17866379686004130, - 64'd2472801959128626, - 64'd341321465710090, - 64'd44117658395661, - 64'd16655495050548274, - 64'd2371002668248148, - 64'd328744863037930, - 64'd43141652534624, - 64'd15495080205241458, - 64'd2270945905806842, - 64'd316291264323041, - 64'd42129783169276, - 64'd14384232414891682, - 64'd2172755029019642, - 64'd303983262307882, - 64'd41087422038183, - 64'd13321990880666632, - 64'd2076539077052086, - 64'd291841332604495, - 64'd40019605208911, - 64'd12307343692121528, - 64'd1982393594214940, - 64'd279883944204480, - 64'd38931045989652}};

	localparam logic signed[63:0] hf[0:1199] = {64'd7838585847808, - 64'd22134781952, - 64'd28777693184, 64'd157109504, 64'd7816469282816, - 64'd66278170624, - 64'd28445626368, 64'd468937216, 64'd7772364603392, - 64'd110045741056, - 64'd27785463808, 64'd773795776, 64'd7706521894912, - 64'd153191858176, - 64'd26804365312, 64'd1067479168, 64'd7619311304704, - 64'd195476406272, - 64'd25512417280, 64'd1346167168, 64'd7511223042048, - 64'd236666617856, - 64'd23922403328, 64'd1606430464, 64'd7382860038144, - 64'd276538851328, - 64'd22049581056, 64'd1845233792, 64'd7234935324672, - 64'd314880131072, - 64'd19911436288, 64'd2059935104, 64'd7068264693760, - 64'd351489753088, - 64'd17527447552, 64'd2248284160, 64'd6883761979392, - 64'd386180317184, - 64'd14918830080, 64'd2408417280, 64'd6682430144512, - 64'd418779267072, - 64'd12108299264, 64'd2538850816, 64'd6465354465280, - 64'd449129578496, - 64'd9119814656, 64'd2638471168, 64'd6233695715328, - 64'd477090775040, - 64'd5978338304, 64'd2706525184, 64'd5988680204288, - 64'd502539649024, - 64'd2709589760, 64'd2742605568, 64'd5731590340608, - 64'd525370720256, 64'd660191040, 64'd2746637568, 64'd5463758340096, - 64'd545496694784, 64'd4104474368, 64'd2718862848, 64'd5186554167296, - 64'd562848792576, 64'd7596666368, 64'd2659820544, 64'd4901378719744, - 64'd577376616448, 64'd11110325248, 64'd2570330112, 64'd4609652293632, - 64'd589048512512, 64'd14619365376, 64'd2451470592, 64'd4312807505920, - 64'd597850980352, 64'd18098251776, 64'd2304559872, 64'd4012278284288, - 64'd603788673024, 64'd21522190336, 64'd2131134208, 64'd3709492264960, - 64'd606883741696, 64'd24867289088, 64'd1932924800, 64'd3405861355520, - 64'd607175639040, 64'd28110718976, 64'd1711836032, 64'd3102774394880, - 64'd604720070656, 64'd31230865408, 64'd1469922944, 64'd2801587453952, - 64'd599588601856, 64'd34207447040, 64'd1209368192, 64'd2503617544192, - 64'd591867478016, 64'd37021638656, 64'd932459648, 64'd2210135015424, - 64'd581657165824, 64'd39656165376, 64'd641567488, 64'd1922356740096, - 64'd569070845952, 64'd42095394816, 64'd339122304, 64'd1641439952896, - 64'd554233692160, 64'd44325408768, 64'd27593422, 64'd1368476221440, - 64'd537281757184, 64'd46334046208, - 64'd290532192, 64'd1104487120896, - 64'd518360662016, 64'd48110952448, - 64'd612770176, 64'd850418991104, - 64'd497624514560, 64'd49647616000, - 64'd936658432, 64'd607139201024, - 64'd475234631680, 64'd50937364480, - 64'd1259775488, 64'd375433035776, - 64'd451358425088, 64'd51975356416, - 64'd1579758208, 64'd156000829440, - 64'd426168025088, 64'd52758601728, - 64'd1894318336, - 64'd50544164864, - 64'd399839166464, 64'd53285892096, - 64'd2201257216, - 64'd243677151232, - 64'd372549812224, 64'd53557784576, - 64'd2498480384, - 64'd422962659328, - 64'd344479170560, 64'd53576552448, - 64'd2784010496, - 64'd588054855680, - 64'd315806285824, 64'd53346115584, - 64'd3055998208, - 64'd738697084928, - 64'd286708989952, 64'd52871962624, - 64'd3312732416, - 64'd874721247232, - 64'd257362853888, 64'd52161089536, - 64'd3552649216, - 64'd996046077952, - 64'd227940040704, 64'd51221897216, - 64'd3774339072, - 64'd1102675443712, - 64'd198608306176, 64'd50064097280, - 64'd3976553216, - 64'd1194695589888, - 64'd169530097664, 64'd48698613760, - 64'd4158207232, - 64'd1272272912384, - 64'd140861603840, 64'd47137476608, - 64'd4318385664, - 64'd1335649501184, - 64'd112752001024, 64'd45393707008, - 64'd4456342528, - 64'd1385140715520, - 64'd85342625792, 64'd43481198592, - 64'd4571503616, - 64'd1421130203136, - 64'd58766360576, 64'd41414606848, - 64'd4663464448, - 64'd1444065837056, - 64'd33147019264, 64'd39209230336, - 64'd4731988992, - 64'd1454455128064, - 64'd8598789120, 64'd36880879616, - 64'd4777006080, - 64'd1452859981824, 64'd14774180864, 64'd34445766656, - 64'd4798607360, - 64'd1439891849216, 64'd36878163968, 64'd31920384000, - 64'd4797039616, - 64'd1416206745600, 64'd57630138368, 64'd29321383936, - 64'd4772701696, - 64'd1382498828288, 64'd76957999104, 64'd26665461760, - 64'd4726133248, - 64'd1339495940096, 64'd94800674816, 64'd23969251328, - 64'd4658012672, - 64'd1287953711104, 64'd111108227072, 64'd21249204224, - 64'd4569144320, - 64'd1228649922560, 64'd125841760256, 64'd18521495552, - 64'd4460450304, - 64'd1162378870784, 64'd138973396992, 64'd15801922560, - 64'd4332963840, - 64'd1089946320896, 64'd150486089728, 64'd13105809408, - 64'd4187813888, - 64'd1012163805184, 64'd160373407744, 64'd10447920128, - 64'd4026220544, - 64'd929843314688, 64'd168639184896, 64'd7842376704, - 64'd3849480192, - 64'd843792711680, 64'd175297282048, 64'd5302585344, - 64'd3658956288, - 64'd754810355712, 64'd180371111936, 64'd2841169920, - 64'd3456067584, - 64'd663680581632, 64'd183893196800, 64'd469909824, - 64'd3242277632, - 64'd571169243136, 64'd185904693248, - 64'd1800311424, - 64'd3019083776, - 64'd478019813376, 64'd186454818816, - 64'd3959552000, - 64'd2788005376, - 64'd384948994048, 64'd185600294912, - 64'd5998848512, - 64'd2550573824, - 64'd292643504128, 64'd183404789760, - 64'd7910247424, - 64'd2308321024, - 64'd201756557312, 64'd179938181120, - 64'd9686825984, - 64'd2062770688, - 64'd112905093120, 64'd175276015616, - 64'd11322705920, - 64'd1815426816, - 64'd26666940416, 64'd169498755072, - 64'd12813063168, - 64'd1567765120, 64'd56421380096, 64'd162691153920, - 64'd14154126336, - 64'd1321224192, 64'd135866646528, 64'd154941538304, - 64'd15343171584, - 64'd1077196544, 64'd211220545536, 64'd146341134336, - 64'd16378506240, - 64'd837020800, 64'd282080968704, 64'd136983355392, - 64'd17259448320, - 64'd601974656, 64'd348092956672, 64'd126963187712, - 64'd17986306048, - 64'd373268192, 64'd408949194752, 64'd116376453120, - 64'd18560339968, - 64'd152037664, 64'd464390422528, 64'd105319194624, - 64'd18983727104, 64'd60659716, 64'd514205384704, 64'd93887053824, - 64'd19259518976, 64'd263850352, 64'd558230274048, 64'd82174640128, - 64'd19391596544, 64'd456648288, 64'd596348305408, 64'd70274949120, - 64'd19384621056, 64'd638258432, 64'd628488667136, 64'd58278825984, - 64'd19243970560, 64'd807979008, 64'd654625341440, 64'd46274449408, - 64'd18975694848, 64'd965203456, 64'd674775564288, 64'd34346823680, - 64'd18586447872, 64'd1109421568, 64'd688998187008, 64'd22577342464, - 64'd18083426304, 64'd1240220032, 64'd697391841280, 64'd11043381248, - 64'd17474308096, 64'd1357281920, 64'd700092710912, - 64'd182086192, - 64'd16767187968, 64'd1460386176, 64'd697272303616, - 64'd11030804480, - 64'd15970506752, 64'd1549406080, 64'd689135026176, - 64'd21439533056, - 64'd15092994048, 64'd1624307200, 64'd675915563008, - 64'd31350288384, - 64'd14143592448, 64'd1685144704, 64'd657876320256, - 64'd40710549504, - 64'd13131402240, 64'd1732060800, 64'd635304542208, - 64'd49473417216, - 64'd12065609728, 64'd1765280128, 64'd608509296640, - 64'd57597730816, - 64'd10955428864, 64'd1785106816, 64'd577819115520, - 64'd65048145920, - 64'd9810040832, 64'd1791919488, 64'd543578456064, - 64'd71795171328, - 64'd8638531584, 64'd1786166784, 64'd506145177600, - 64'd77815152640, - 64'd7449839616, 64'd1768361856, 64'd465887559680, - 64'd83090268160, - 64'd6252702208, 64'd1739077632, 64'd423181254656, - 64'd87608377344, - 64'd5055602176, 64'd1698940800, 64'd378406633472, - 64'd91362983936, - 64'd3866723584, 64'd1648625920, 64'd331945902080, - 64'd94353039360, - 64'd2693908224, 64'd1588849920, 64'd284180545536, - 64'd96582770688, - 64'd1544613632, 64'd1520366336, 64'd235488575488, - 64'd98061484032, - 64'd425878816, 64'd1443958144, 64'd186242170880, - 64'd98803326976, 64'd655708864, 64'd1360433152, 64'd136805277696, - 64'd98827001856, 64'd1694041216, 64'd1270616832, 64'd87531372544, - 64'd98155536384, 64'd2683514112, 64'd1175347072, 64'd38761455616, - 64'd96815923200, 64'd3619046400, 64'd1075467904, - 64'd9177933824, - 64'd94838857728, 64'd4496097280, 64'd971824320, - 64'd55976439808, - 64'd92258361344, 64'd5310675968, 64'd865255936, - 64'd101341495296, - 64'd89111461888, 64'd6059353088, 64'd756592576, - 64'd144999710720, - 64'd85437849600, 64'd6739259392, 64'd646648640, - 64'd186698153984, - 64'd81279500288, 64'd7348090880, 64'd536218368, - 64'd226205335552, - 64'd76680314880, 64'd7884102144, 64'd426071456, - 64'd263312162816, - 64'd71685799936, 64'd8346099200, 64'd316948736, - 64'd297832611840, - 64'd66342629376, 64'd8733430784, 64'd209558320, - 64'd329604202496, - 64'd60698370048, 64'd9045970944, 64'd104572016, - 64'd358488408064, - 64'd54801076224, 64'd9284107264, 64'd2622117, - 64'd384370769920, - 64'd48698970112, 64'd9448714240, - 64'd95701408, - 64'd407160881152, - 64'd42440110080, 64'd9541138432, - 64'd189853392, - 64'd426792321024, - 64'd36072067072, 64'd9563166720, - 64'd279335552, - 64'd443222228992, - 64'd29641613312, 64'd9517003776, - 64'd363698272, - 64'd456430845952, - 64'd23194449920, 64'd9405243392, - 64'd442541760, - 64'd466420989952, - 64'd16774914048, 64'd9230835712, - 64'd515517248, - 64'd473217204224, - 64'd10425733120, 64'd8997056512, - 64'd582327424, - 64'd476865003520, - 64'd4187790080, 64'd8707474432, - 64'd642726784, - 64'd477429760000, 64'd1900096640, 64'd8365917696, - 64'd696521408, - 64'd474995785728, 64'd7801364992, 64'd7976438784, - 64'd743568576, - 64'd469664989184, 64'd13481884672, 64'd7543281152, - 64'd783776000, - 64'd461555793920, 64'd18910107648, 64'd7070841856, - 64'd817100608, - 64'd450801598464, 64'd24057192448, 64'd6563639808, - 64'd843547520, - 64'd437549662208, 64'd28897122304, 64'd6026279936, - 64'd863167872, - 64'd421959434240, 64'd33406773248, 64'd5463418880, - 64'd876057536, - 64'd404201209856, 64'd37565992960, 64'd4879733248, - 64'd882354496, - 64'd384454656000, 64'd41357627392, 64'd4279885568, - 64'd882236544, - 64'd362907205632, 64'd44767539200, 64'd3668495872, - 64'd875919168, - 64'd339752583168, 64'd47784624128, 64'd3050110720, - 64'd863652352, - 64'd315189428224, 64'd50400759808, 64'd2429174528, - 64'd845718144, - 64'd289419558912, 64'd52610781184, 64'd1810003712, - 64'd822427328, - 64'd262646759424, 64'd54412427264, 64'd1196761984, - 64'd794116736, - 64'd235075190784, 64'd55806234624, 64'd593437184, - 64'd761145856, - 64'd206908047360, 64'd56795480064, 64'd3820039, - 64'd723893696, - 64'd178346278912, 64'd57386037248, - 64'd568514688, - 64'd682755840, - 64'd149587197952, 64'd57586274304, - 64'd1120225152, - 64'd638140992, - 64'd120823414784, 64'd57406910464, - 64'd1648217344, - 64'd590467712, - 64'd92241559552, 64'd56860872704, - 64'd2149657600, - 64'd540161664, - 64'd64021319680, 64'd55963131904, - 64'd2621983744, - 64'd487652064, - 64'd36334411776, 64'd54730534912, - 64'd3062912256, - 64'd433369056, - 64'd9343685632, 64'd53181644800, - 64'd3470446080, - 64'd377740576, 64'd16797673472, 64'd51336544256, - 64'd3842877184, - 64'd321189600, 64'd41946865664, 64'd49216663552, - 64'd4178790144, - 64'd264131488, 64'd65972105216, 64'd46844592128, - 64'd4477060608, - 64'd206971392, 64'd88753152000, 64'd44243890176, - 64'd4736854016, - 64'd150101952, 64'd110181744640, 64'd41438887936, - 64'd4957623296, - 64'd93900968, 64'd130161942528, 64'd38454513664, - 64'd5139099648, - 64'd38729428, 64'd148610383872, 64'd35316113408, - 64'd5281288704, 64'd15070397, 64'd165456445440, 64'd32049231872, - 64'd5384460800, 64'd67176656, 64'd180642283520, 64'd28679483392, - 64'd5449138176, 64'd117289376, 64'd194122842112, 64'd25232340992, - 64'd5476087296, 64'd165131808, 64'd205865746432, 64'd21732986880, - 64'd5466302464, 64'd210451488, 64'd215851089920, 64'd18206152704, - 64'd5420994048, 64'd253021136, 64'd224071172096, 64'd14675965952, - 64'd5341570560, 64'd292639424, 64'd230530236416, 64'd11165807616, - 64'd5229625856, 64'd329131392, 64'd235243929600, 64'd7698181120, - 64'd5086921728, 64'd362348864, 64'd238238957568, 64'd4294591744, - 64'd4915367936, 64'd392170432, 64'd239552479232, 64'd975431552, - 64'd4717009408, 64'd418501568, 64'd239231549440, - 64'd2240118784, - 64'd4494003712, 64'd441274240, 64'd237332512768, - 64'd5334179840, - 64'd4248604672, 64'd460446592, 64'd233920282624, - 64'd8290250240, - 64'd3983145216, 64'd476002368, 64'd229067702272, - 64'd11093274624, - 64'd3700017920, 64'd487950112, 64'd222854709248, - 64'd13729694720, - 64'd3401656832, 64'd496322432, 64'd215367729152, - 64'd16187494400, - 64'd3090520832, 64'd501174912, 64'd206698692608, - 64'd18456229888, - 64'd2769075712, 64'd502584992, 64'd196944461824, - 64'd20527046656, - 64'd2439777280, 64'd500650752, 64'd186205831168, - 64'd22392690688, - 64'd2105056128, 64'd495489664, 64'd174586904576, - 64'd24047501312, - 64'd1767301120, 64'd487237024, 64'd162194161664, - 64'd25487403008, - 64'd1428845312, 64'd476044576, 64'd149135753216, - 64'd26709876736, - 64'd1091952000, 64'd462079008, 64'd135520722944, - 64'd27713929216, - 64'd758801984, 64'd445520128, 64'd121458196480, - 64'd28500049920, - 64'd431481408, 64'd426559552, 64'd107056726016, - 64'd29070161920, - 64'd111970936, 64'd405398752, 64'd92423544832, - 64'd29427556352, 64'd197864096, 64'd382247584, 64'd77663920128, - 64'd29576835072, 64'd496282400, 64'd357322464, 64'd62880497664, - 64'd29523832832, 64'd781674496, 64'd330844800, 64'd48172716032, - 64'd29275539456, 64'd1052569088, 64'd303039392, 64'd33636249600, - 64'd28840015872, 64'd1307638528, 64'd274132608, 64'd19362488320, - 64'd28226306048, 64'd1545703040, 64'd244351072, 64'd5438078976, - 64'd27444344832, 64'd1765733888, 64'd213919968, - 64'd8055504896, - 64'd26504861696, 64'd1966855424, 64'd183061680, - 64'd21042335744, - 64'd25419290624, 64'd2148345856, 64'd151994288, - 64'd33452351488, - 64'd24199659520, 64'd2309637120, 64'd120930336, - 64'd45221638144, - 64'd22858500096, 64'd2450314240, 64'd90075568, - 64'd56292646912, - 64'd21408743424, 64'd2570112000, 64'd59627728, - 64'd66614386688, - 64'd19863625728, 64'd2668913152, 64'd29775562, - 64'd76142518272, - 64'd18236581888, 64'd2746743552, 64'd697786, - 64'd84839473152, - 64'd16541160448, 64'd2803768576, - 64'd27437750, - 64'd92674449408, - 64'd14790919168, 64'd2840285696, - 64'd54474848, - 64'd99623403520, - 64'd12999341056, 64'd2856719616, - 64'd80269632, - 64'd105669025792, - 64'd11179744256, 64'd2853614848, - 64'd104691112, - 64'd110800576512, - 64'd9345202176, 64'd2831628544, - 64'd127621640, - 64'd115013779456, - 64'd7508456960, 64'd2791522048, - 64'd148957264, - 64'd118310641664, - 64'd5681853440, 64'd2734152704, - 64'd168607984, - 64'd120699232256, - 64'd3877264384, 64'd2660464896, - 64'd186497920, - 64'd122193403904, - 64'd2106029312, 64'd2571481344, - 64'd202565360, - 64'd122812547072, - 64'd378894784, 64'd2468293376, - 64'd216762656, - 64'd122581278720, 64'd1294037120, 64'd2352050944, - 64'd229056208, - 64'd121529065472, 64'd2903355648, 64'd2223954432, - 64'd239426112, - 64'd119689928704, 64'd4440381440, 64'd2085244032, - 64'd247865936, - 64'd117102018560, 64'd5897201664, 64'd1937189760, - 64'd254382288, - 64'd113807253504, 64'd7266695168, 64'd1781083520, - 64'd258994368, - 64'd109850902528, 64'd8542557696, 64'd1618228224, - 64'd261733440, - 64'd105281200128, 64'd9719314432, 64'd1449929984, - 64'd262642192, - 64'd100148871168, 64'd10792333312, 64'd1277488256, - 64'd261774160, - 64'd94506778624, 64'd11757822976, 64'd1102188160, - 64'd259192944, - 64'd88409464832, 64'd12612836352, 64'd925292096, - 64'd254971488, - 64'd81912717312, 64'd13355259904, 64'd748031936, - 64'd249191312, - 64'd75073200128, 64'd13983799296, 64'd571602112, - 64'd241941664, - 64'd67947999232, 64'd14497965056, 64'd397152512, - 64'd233318704, - 64'd60594270208, 64'd14898048000, 64'd225782496, - 64'd223424592, - 64'd53068820480, 64'd15185090560, 64'd58535152, - 64'd212366656, - 64'd45427761152, 64'd15360858112, - 64'd103607888, - 64'd200256496, - 64'd37726138368, 64'd15427800064, - 64'd259730960, - 64'd187209104, - 64'd30017622016, 64'd15389016064, - 64'd408988352, - 64'd173341968, - 64'd22354171904, 64'd15248207872, - 64'd550607616, - 64'd158774256, - 64'd14785753088, 64'd15009643520, - 64'd683892544, - 64'd143625904, - 64'd7360073728, 64'd14678099968, - 64'd808224960, - 64'd128016848, - 64'd122326760, 64'd14258824192, - 64'd923066752, - 64'd112066168, 64'd6885020160, 64'd13757478912, - 64'd1027960576, - 64'd95891384, 64'd13622423552, 64'd13180087296, - 64'd1122530432, - 64'd79607672, 64'd20053434368, 64'd12532989952, - 64'd1206481152, - 64'd63327192, 64'd26144839680, 64'd11822783488, - 64'd1279598592, - 64'd47158456, 64'd31866779648, 64'd11056274432, - 64'd1341747456, - 64'd31205682, 64'd37192835072, 64'd10240421888, - 64'd1392870272, - 64'd15568271, 64'd42100101120, 64'd9382290432, - 64'd1432985088, - 64'd340284, 64'd46569213952, 64'd8488998400, - 64'd1462182656, 64'd14390004, 64'd50584375296, 64'd7567664640, - 64'd1480623872, 64'd28540510, 64'd54133334016, 64'd6625367552, - 64'd1488536064, 64'd42035688, 64'd57207365632, 64'd5669093376, - 64'd1486209792, 64'd54806824, 64'd59801194496, 64'd4705696256, - 64'd1473994240, 64'd66792264, 64'd61912944640, 64'd3741853952, - 64'd1452293376, 64'd77937600, 64'd63544012800, 64'd2784031744, - 64'd1421561344, 64'd88195824, 64'd64698974208, 64'd1838443904, - 64'd1382297856, 64'd97527336, 64'd65385447424, 64'd911020864, - 64'd1335043584, 64'd105900048, 64'd65613926400, 64'd7379710, - 64'd1280374656, 64'd113289296, 64'd65397641216, - 64'd867204224, - 64'd1218898048, 64'd119677792, 64'd64752361472, - 64'd1707821056, - 64'd1151246848, 64'd125055480, 64'd63696216064, - 64'd2509947136, - 64'd1078074240, 64'd129419384, 64'd62249496576, - 64'd3269463296, - 64'd1000049600, 64'd132773400, 64'd60434452480, - 64'd3982668544, - 64'd917852672, 64'd135128032, 64'd58275078144, - 64'd4646291968, - 64'd832168896, 64'd136500128, 64'd55796891648, - 64'd5257499648, - 64'd743684992, 64'd136912544, 64'd53026709504, - 64'd5813900800, - 64'd653083904, 64'd136393792, 64'd49992445952, - 64'd6313548288, - 64'd561040576, 64'd134977664, 64'd46722871296, - 64'd6754936320, - 64'd468217632, 64'd132702888, 64'd43247403008, - 64'd7136999424, - 64'd375261408, 64'd129612640, 64'd39595872256, - 64'd7459101696, - 64'd282798048, 64'd125754136, 64'd35798339584, - 64'd7721029120, - 64'd191430208, 64'd121178200, 64'd31884855296, - 64'd7922977280, - 64'd101733480, 64'd115938792, 64'd27885277184, - 64'd8065535488, - 64'd14253701, 64'd110092552, 64'd23829073920, - 64'd8149671936, 64'd70495888, 64'd103698320, 64'd19745140736, - 64'd8176712704, 64'd152036944, 64'd96816696, 64'd15661621248, - 64'd8148323328, 64'd229928128, 64'd89509568, 64'd11605748736, - 64'd8066485760, 64'd303766784, 64'd81839656, 64'd7603688960, - 64'd7933474816, 64'd373190432, 64'd73870048, 64'd3680404224, - 64'd7751833600, 64'd437877920, 64'd65663800, - 64'd140476864, - 64'd7524347392, 64'd497550080, 64'd57283504, - 64'd3836774656, - 64'd7254018048, 64'd551970432, 64'd48790868, - 64'd7387857920, - 64'd6944036352, 64'd600945152, 64'd40246348, - 64'd10774731776, - 64'd6597754880, 64'd644323200, 64'd31708794, - 64'd13980114944, - 64'd6218660352, 64'd681995840, 64'd23235080, - 64'd16988492800, - 64'd5810344448, 64'd713896000, 64'd14879819, - 64'd19786172416, - 64'd5376479744, 64'd739997248, 64'd6695052, - 64'd22361307136, - 64'd4920788992, 64'd760312896, - 64'd1270005, - 64'd24703920128, - 64'd4447020544, 64'd774894464, - 64'd8969208, - 64'd26805911552, - 64'd3958922496, 64'd783830144, - 64'd16359686, - 64'd28661049344, - 64'd3460217344, 64'd787242880, - 64'd23402022, - 64'd30264948736, - 64'd2954577408, 64'd785288704, - 64'd30060408, - 64'd31615045632, - 64'd2445602560, 64'd778154368, - 64'd36302760, - 64'd32710555648, - 64'd1936798720, 64'd766055168, - 64'd42100824, - 64'd33552416768, - 64'd1431556480, 64'd749232704, - 64'd47430228, - 64'd34143229952, - 64'd933133504, 64'd727952128, - 64'd52270520, - 64'd34487185408, - 64'd444635872, 64'd702499968, - 64'd56605188, - 64'd34589990912, 64'd30996946, 64'd673181248, - 64'd60421624, - 64'd34458779648, 64'd491006656, 64'd640316992, - 64'd63711108, - 64'd34102003712, 64'd932828672, 64'd604241408, - 64'd66468712, - 64'd33529362432, 64'd1354102784, 64'd565299456, - 64'd68693224, - 64'd32751673344, 64'd1752682880, 64'd523844032, - 64'd70387048, - 64'd31780775936, 64'd2126643328, 64'd480233312, - 64'd71556032, - 64'd30629410816, 64'd2474285568, 64'd434828384, - 64'd72209368, - 64'd29311117312, 64'd2794141952, 64'd387990528, - 64'd72359368, - 64'd27840104448, 64'd3084977920, 64'd340078944, - 64'd72021344, - 64'd26231142400, 64'd3345792256, 64'd291448352, - 64'd71213336, - 64'd24499443712, 64'd3575817216, 64'd242446768, - 64'd69955968, - 64'd22660548608, 64'd3774514944, 64'd193413440, - 64'd68272184, - 64'd20730206208, 64'd3941574912, 64'd144676800, - 64'd66187028, - 64'd18724265984, 64'd4076907264, 64'd96552704, - 64'd63727432, - 64'd16658572288, 64'd4180636928, 64'd49342632, - 64'd60921944, - 64'd14548849664, 64'd4253096448, 64'd3332228, - 64'd57800504, - 64'd12410608640, 64'd4294816000, - 64'd41210148, - 64'd54394188, - 64'd10259047424, 64'd4306513408, - 64'd84034640, - 64'd50734972, - 64'd8108961280, 64'd4289084160, - 64'd124910944, - 64'd46855484, - 64'd5974653440, 64'd4243589120, - 64'd163629248, - 64'd42788764};

	localparam logic signed[63:0] hb[0:1199] = {64'd7838585847808, 64'd22134781952, - 64'd28777693184, - 64'd157109504, 64'd7816469282816, 64'd66278170624, - 64'd28445626368, - 64'd468937216, 64'd7772364603392, 64'd110045741056, - 64'd27785463808, - 64'd773795776, 64'd7706521894912, 64'd153191858176, - 64'd26804365312, - 64'd1067479168, 64'd7619311304704, 64'd195476406272, - 64'd25512417280, - 64'd1346167168, 64'd7511223042048, 64'd236666617856, - 64'd23922403328, - 64'd1606430464, 64'd7382860038144, 64'd276538851328, - 64'd22049581056, - 64'd1845233792, 64'd7234935324672, 64'd314880131072, - 64'd19911436288, - 64'd2059935104, 64'd7068264693760, 64'd351489753088, - 64'd17527447552, - 64'd2248284160, 64'd6883761979392, 64'd386180317184, - 64'd14918830080, - 64'd2408417280, 64'd6682430144512, 64'd418779267072, - 64'd12108299264, - 64'd2538850816, 64'd6465354465280, 64'd449129578496, - 64'd9119814656, - 64'd2638471168, 64'd6233695715328, 64'd477090775040, - 64'd5978338304, - 64'd2706525184, 64'd5988680204288, 64'd502539649024, - 64'd2709589760, - 64'd2742605568, 64'd5731590340608, 64'd525370720256, 64'd660191040, - 64'd2746637568, 64'd5463758340096, 64'd545496694784, 64'd4104474368, - 64'd2718862848, 64'd5186554167296, 64'd562848792576, 64'd7596666368, - 64'd2659820544, 64'd4901378719744, 64'd577376616448, 64'd11110325248, - 64'd2570330112, 64'd4609652293632, 64'd589048512512, 64'd14619365376, - 64'd2451470592, 64'd4312807505920, 64'd597850980352, 64'd18098251776, - 64'd2304559872, 64'd4012278284288, 64'd603788673024, 64'd21522190336, - 64'd2131134208, 64'd3709492264960, 64'd606883741696, 64'd24867289088, - 64'd1932924800, 64'd3405861355520, 64'd607175639040, 64'd28110718976, - 64'd1711836032, 64'd3102774394880, 64'd604720070656, 64'd31230865408, - 64'd1469922944, 64'd2801587453952, 64'd599588601856, 64'd34207447040, - 64'd1209368192, 64'd2503617544192, 64'd591867478016, 64'd37021638656, - 64'd932459648, 64'd2210135015424, 64'd581657165824, 64'd39656165376, - 64'd641567488, 64'd1922356740096, 64'd569070845952, 64'd42095394816, - 64'd339122304, 64'd1641439952896, 64'd554233692160, 64'd44325408768, - 64'd27593422, 64'd1368476221440, 64'd537281757184, 64'd46334046208, 64'd290532192, 64'd1104487120896, 64'd518360662016, 64'd48110952448, 64'd612770176, 64'd850418991104, 64'd497624514560, 64'd49647616000, 64'd936658432, 64'd607139201024, 64'd475234631680, 64'd50937364480, 64'd1259775488, 64'd375433035776, 64'd451358425088, 64'd51975356416, 64'd1579758208, 64'd156000829440, 64'd426168025088, 64'd52758601728, 64'd1894318336, - 64'd50544164864, 64'd399839166464, 64'd53285892096, 64'd2201257216, - 64'd243677151232, 64'd372549812224, 64'd53557784576, 64'd2498480384, - 64'd422962659328, 64'd344479170560, 64'd53576552448, 64'd2784010496, - 64'd588054855680, 64'd315806285824, 64'd53346115584, 64'd3055998208, - 64'd738697084928, 64'd286708989952, 64'd52871962624, 64'd3312732416, - 64'd874721247232, 64'd257362853888, 64'd52161089536, 64'd3552649216, - 64'd996046077952, 64'd227940040704, 64'd51221897216, 64'd3774339072, - 64'd1102675443712, 64'd198608306176, 64'd50064097280, 64'd3976553216, - 64'd1194695589888, 64'd169530097664, 64'd48698613760, 64'd4158207232, - 64'd1272272912384, 64'd140861603840, 64'd47137476608, 64'd4318385664, - 64'd1335649501184, 64'd112752001024, 64'd45393707008, 64'd4456342528, - 64'd1385140715520, 64'd85342625792, 64'd43481198592, 64'd4571503616, - 64'd1421130203136, 64'd58766360576, 64'd41414606848, 64'd4663464448, - 64'd1444065837056, 64'd33147019264, 64'd39209230336, 64'd4731988992, - 64'd1454455128064, 64'd8598789120, 64'd36880879616, 64'd4777006080, - 64'd1452859981824, - 64'd14774180864, 64'd34445766656, 64'd4798607360, - 64'd1439891849216, - 64'd36878163968, 64'd31920384000, 64'd4797039616, - 64'd1416206745600, - 64'd57630138368, 64'd29321383936, 64'd4772701696, - 64'd1382498828288, - 64'd76957999104, 64'd26665461760, 64'd4726133248, - 64'd1339495940096, - 64'd94800674816, 64'd23969251328, 64'd4658012672, - 64'd1287953711104, - 64'd111108227072, 64'd21249204224, 64'd4569144320, - 64'd1228649922560, - 64'd125841760256, 64'd18521495552, 64'd4460450304, - 64'd1162378870784, - 64'd138973396992, 64'd15801922560, 64'd4332963840, - 64'd1089946320896, - 64'd150486089728, 64'd13105809408, 64'd4187813888, - 64'd1012163805184, - 64'd160373407744, 64'd10447920128, 64'd4026220544, - 64'd929843314688, - 64'd168639184896, 64'd7842376704, 64'd3849480192, - 64'd843792711680, - 64'd175297282048, 64'd5302585344, 64'd3658956288, - 64'd754810355712, - 64'd180371111936, 64'd2841169920, 64'd3456067584, - 64'd663680581632, - 64'd183893196800, 64'd469909824, 64'd3242277632, - 64'd571169243136, - 64'd185904693248, - 64'd1800311424, 64'd3019083776, - 64'd478019813376, - 64'd186454818816, - 64'd3959552000, 64'd2788005376, - 64'd384948994048, - 64'd185600294912, - 64'd5998848512, 64'd2550573824, - 64'd292643504128, - 64'd183404789760, - 64'd7910247424, 64'd2308321024, - 64'd201756557312, - 64'd179938181120, - 64'd9686825984, 64'd2062770688, - 64'd112905093120, - 64'd175276015616, - 64'd11322705920, 64'd1815426816, - 64'd26666940416, - 64'd169498755072, - 64'd12813063168, 64'd1567765120, 64'd56421380096, - 64'd162691153920, - 64'd14154126336, 64'd1321224192, 64'd135866646528, - 64'd154941538304, - 64'd15343171584, 64'd1077196544, 64'd211220545536, - 64'd146341134336, - 64'd16378506240, 64'd837020800, 64'd282080968704, - 64'd136983355392, - 64'd17259448320, 64'd601974656, 64'd348092956672, - 64'd126963187712, - 64'd17986306048, 64'd373268192, 64'd408949194752, - 64'd116376453120, - 64'd18560339968, 64'd152037664, 64'd464390422528, - 64'd105319194624, - 64'd18983727104, - 64'd60659716, 64'd514205384704, - 64'd93887053824, - 64'd19259518976, - 64'd263850352, 64'd558230274048, - 64'd82174640128, - 64'd19391596544, - 64'd456648288, 64'd596348305408, - 64'd70274949120, - 64'd19384621056, - 64'd638258432, 64'd628488667136, - 64'd58278825984, - 64'd19243970560, - 64'd807979008, 64'd654625341440, - 64'd46274449408, - 64'd18975694848, - 64'd965203456, 64'd674775564288, - 64'd34346823680, - 64'd18586447872, - 64'd1109421568, 64'd688998187008, - 64'd22577342464, - 64'd18083426304, - 64'd1240220032, 64'd697391841280, - 64'd11043381248, - 64'd17474308096, - 64'd1357281920, 64'd700092710912, 64'd182086192, - 64'd16767187968, - 64'd1460386176, 64'd697272303616, 64'd11030804480, - 64'd15970506752, - 64'd1549406080, 64'd689135026176, 64'd21439533056, - 64'd15092994048, - 64'd1624307200, 64'd675915563008, 64'd31350288384, - 64'd14143592448, - 64'd1685144704, 64'd657876320256, 64'd40710549504, - 64'd13131402240, - 64'd1732060800, 64'd635304542208, 64'd49473417216, - 64'd12065609728, - 64'd1765280128, 64'd608509296640, 64'd57597730816, - 64'd10955428864, - 64'd1785106816, 64'd577819115520, 64'd65048145920, - 64'd9810040832, - 64'd1791919488, 64'd543578456064, 64'd71795171328, - 64'd8638531584, - 64'd1786166784, 64'd506145177600, 64'd77815152640, - 64'd7449839616, - 64'd1768361856, 64'd465887559680, 64'd83090268160, - 64'd6252702208, - 64'd1739077632, 64'd423181254656, 64'd87608377344, - 64'd5055602176, - 64'd1698940800, 64'd378406633472, 64'd91362983936, - 64'd3866723584, - 64'd1648625920, 64'd331945902080, 64'd94353039360, - 64'd2693908224, - 64'd1588849920, 64'd284180545536, 64'd96582770688, - 64'd1544613632, - 64'd1520366336, 64'd235488575488, 64'd98061484032, - 64'd425878816, - 64'd1443958144, 64'd186242170880, 64'd98803326976, 64'd655708864, - 64'd1360433152, 64'd136805277696, 64'd98827001856, 64'd1694041216, - 64'd1270616832, 64'd87531372544, 64'd98155536384, 64'd2683514112, - 64'd1175347072, 64'd38761455616, 64'd96815923200, 64'd3619046400, - 64'd1075467904, - 64'd9177933824, 64'd94838857728, 64'd4496097280, - 64'd971824320, - 64'd55976439808, 64'd92258361344, 64'd5310675968, - 64'd865255936, - 64'd101341495296, 64'd89111461888, 64'd6059353088, - 64'd756592576, - 64'd144999710720, 64'd85437849600, 64'd6739259392, - 64'd646648640, - 64'd186698153984, 64'd81279500288, 64'd7348090880, - 64'd536218368, - 64'd226205335552, 64'd76680314880, 64'd7884102144, - 64'd426071456, - 64'd263312162816, 64'd71685799936, 64'd8346099200, - 64'd316948736, - 64'd297832611840, 64'd66342629376, 64'd8733430784, - 64'd209558320, - 64'd329604202496, 64'd60698370048, 64'd9045970944, - 64'd104572016, - 64'd358488408064, 64'd54801076224, 64'd9284107264, - 64'd2622117, - 64'd384370769920, 64'd48698970112, 64'd9448714240, 64'd95701408, - 64'd407160881152, 64'd42440110080, 64'd9541138432, 64'd189853392, - 64'd426792321024, 64'd36072067072, 64'd9563166720, 64'd279335552, - 64'd443222228992, 64'd29641613312, 64'd9517003776, 64'd363698272, - 64'd456430845952, 64'd23194449920, 64'd9405243392, 64'd442541760, - 64'd466420989952, 64'd16774914048, 64'd9230835712, 64'd515517248, - 64'd473217204224, 64'd10425733120, 64'd8997056512, 64'd582327424, - 64'd476865003520, 64'd4187790080, 64'd8707474432, 64'd642726784, - 64'd477429760000, - 64'd1900096640, 64'd8365917696, 64'd696521408, - 64'd474995785728, - 64'd7801364992, 64'd7976438784, 64'd743568576, - 64'd469664989184, - 64'd13481884672, 64'd7543281152, 64'd783776000, - 64'd461555793920, - 64'd18910107648, 64'd7070841856, 64'd817100608, - 64'd450801598464, - 64'd24057192448, 64'd6563639808, 64'd843547520, - 64'd437549662208, - 64'd28897122304, 64'd6026279936, 64'd863167872, - 64'd421959434240, - 64'd33406773248, 64'd5463418880, 64'd876057536, - 64'd404201209856, - 64'd37565992960, 64'd4879733248, 64'd882354496, - 64'd384454656000, - 64'd41357627392, 64'd4279885568, 64'd882236544, - 64'd362907205632, - 64'd44767539200, 64'd3668495872, 64'd875919168, - 64'd339752583168, - 64'd47784624128, 64'd3050110720, 64'd863652352, - 64'd315189428224, - 64'd50400759808, 64'd2429174528, 64'd845718144, - 64'd289419558912, - 64'd52610781184, 64'd1810003712, 64'd822427328, - 64'd262646759424, - 64'd54412427264, 64'd1196761984, 64'd794116736, - 64'd235075190784, - 64'd55806234624, 64'd593437184, 64'd761145856, - 64'd206908047360, - 64'd56795480064, 64'd3820039, 64'd723893696, - 64'd178346278912, - 64'd57386037248, - 64'd568514688, 64'd682755840, - 64'd149587197952, - 64'd57586274304, - 64'd1120225152, 64'd638140992, - 64'd120823414784, - 64'd57406910464, - 64'd1648217344, 64'd590467712, - 64'd92241559552, - 64'd56860872704, - 64'd2149657600, 64'd540161664, - 64'd64021319680, - 64'd55963131904, - 64'd2621983744, 64'd487652064, - 64'd36334411776, - 64'd54730534912, - 64'd3062912256, 64'd433369056, - 64'd9343685632, - 64'd53181644800, - 64'd3470446080, 64'd377740576, 64'd16797673472, - 64'd51336544256, - 64'd3842877184, 64'd321189600, 64'd41946865664, - 64'd49216663552, - 64'd4178790144, 64'd264131488, 64'd65972105216, - 64'd46844592128, - 64'd4477060608, 64'd206971392, 64'd88753152000, - 64'd44243890176, - 64'd4736854016, 64'd150101952, 64'd110181744640, - 64'd41438887936, - 64'd4957623296, 64'd93900968, 64'd130161942528, - 64'd38454513664, - 64'd5139099648, 64'd38729428, 64'd148610383872, - 64'd35316113408, - 64'd5281288704, - 64'd15070397, 64'd165456445440, - 64'd32049231872, - 64'd5384460800, - 64'd67176656, 64'd180642283520, - 64'd28679483392, - 64'd5449138176, - 64'd117289376, 64'd194122842112, - 64'd25232340992, - 64'd5476087296, - 64'd165131808, 64'd205865746432, - 64'd21732986880, - 64'd5466302464, - 64'd210451488, 64'd215851089920, - 64'd18206152704, - 64'd5420994048, - 64'd253021136, 64'd224071172096, - 64'd14675965952, - 64'd5341570560, - 64'd292639424, 64'd230530236416, - 64'd11165807616, - 64'd5229625856, - 64'd329131392, 64'd235243929600, - 64'd7698181120, - 64'd5086921728, - 64'd362348864, 64'd238238957568, - 64'd4294591744, - 64'd4915367936, - 64'd392170432, 64'd239552479232, - 64'd975431552, - 64'd4717009408, - 64'd418501568, 64'd239231549440, 64'd2240118784, - 64'd4494003712, - 64'd441274240, 64'd237332512768, 64'd5334179840, - 64'd4248604672, - 64'd460446592, 64'd233920282624, 64'd8290250240, - 64'd3983145216, - 64'd476002368, 64'd229067702272, 64'd11093274624, - 64'd3700017920, - 64'd487950112, 64'd222854709248, 64'd13729694720, - 64'd3401656832, - 64'd496322432, 64'd215367729152, 64'd16187494400, - 64'd3090520832, - 64'd501174912, 64'd206698692608, 64'd18456229888, - 64'd2769075712, - 64'd502584992, 64'd196944461824, 64'd20527046656, - 64'd2439777280, - 64'd500650752, 64'd186205831168, 64'd22392690688, - 64'd2105056128, - 64'd495489664, 64'd174586904576, 64'd24047501312, - 64'd1767301120, - 64'd487237024, 64'd162194161664, 64'd25487403008, - 64'd1428845312, - 64'd476044576, 64'd149135753216, 64'd26709876736, - 64'd1091952000, - 64'd462079008, 64'd135520722944, 64'd27713929216, - 64'd758801984, - 64'd445520128, 64'd121458196480, 64'd28500049920, - 64'd431481408, - 64'd426559552, 64'd107056726016, 64'd29070161920, - 64'd111970936, - 64'd405398752, 64'd92423544832, 64'd29427556352, 64'd197864096, - 64'd382247584, 64'd77663920128, 64'd29576835072, 64'd496282400, - 64'd357322464, 64'd62880497664, 64'd29523832832, 64'd781674496, - 64'd330844800, 64'd48172716032, 64'd29275539456, 64'd1052569088, - 64'd303039392, 64'd33636249600, 64'd28840015872, 64'd1307638528, - 64'd274132608, 64'd19362488320, 64'd28226306048, 64'd1545703040, - 64'd244351072, 64'd5438078976, 64'd27444344832, 64'd1765733888, - 64'd213919968, - 64'd8055504896, 64'd26504861696, 64'd1966855424, - 64'd183061680, - 64'd21042335744, 64'd25419290624, 64'd2148345856, - 64'd151994288, - 64'd33452351488, 64'd24199659520, 64'd2309637120, - 64'd120930336, - 64'd45221638144, 64'd22858500096, 64'd2450314240, - 64'd90075568, - 64'd56292646912, 64'd21408743424, 64'd2570112000, - 64'd59627728, - 64'd66614386688, 64'd19863625728, 64'd2668913152, - 64'd29775562, - 64'd76142518272, 64'd18236581888, 64'd2746743552, - 64'd697786, - 64'd84839473152, 64'd16541160448, 64'd2803768576, 64'd27437750, - 64'd92674449408, 64'd14790919168, 64'd2840285696, 64'd54474848, - 64'd99623403520, 64'd12999341056, 64'd2856719616, 64'd80269632, - 64'd105669025792, 64'd11179744256, 64'd2853614848, 64'd104691112, - 64'd110800576512, 64'd9345202176, 64'd2831628544, 64'd127621640, - 64'd115013779456, 64'd7508456960, 64'd2791522048, 64'd148957264, - 64'd118310641664, 64'd5681853440, 64'd2734152704, 64'd168607984, - 64'd120699232256, 64'd3877264384, 64'd2660464896, 64'd186497920, - 64'd122193403904, 64'd2106029312, 64'd2571481344, 64'd202565360, - 64'd122812547072, 64'd378894784, 64'd2468293376, 64'd216762656, - 64'd122581278720, - 64'd1294037120, 64'd2352050944, 64'd229056208, - 64'd121529065472, - 64'd2903355648, 64'd2223954432, 64'd239426112, - 64'd119689928704, - 64'd4440381440, 64'd2085244032, 64'd247865936, - 64'd117102018560, - 64'd5897201664, 64'd1937189760, 64'd254382288, - 64'd113807253504, - 64'd7266695168, 64'd1781083520, 64'd258994368, - 64'd109850902528, - 64'd8542557696, 64'd1618228224, 64'd261733440, - 64'd105281200128, - 64'd9719314432, 64'd1449929984, 64'd262642192, - 64'd100148871168, - 64'd10792333312, 64'd1277488256, 64'd261774160, - 64'd94506778624, - 64'd11757822976, 64'd1102188160, 64'd259192944, - 64'd88409464832, - 64'd12612836352, 64'd925292096, 64'd254971488, - 64'd81912717312, - 64'd13355259904, 64'd748031936, 64'd249191312, - 64'd75073200128, - 64'd13983799296, 64'd571602112, 64'd241941664, - 64'd67947999232, - 64'd14497965056, 64'd397152512, 64'd233318704, - 64'd60594270208, - 64'd14898048000, 64'd225782496, 64'd223424592, - 64'd53068820480, - 64'd15185090560, 64'd58535152, 64'd212366656, - 64'd45427761152, - 64'd15360858112, - 64'd103607888, 64'd200256496, - 64'd37726138368, - 64'd15427800064, - 64'd259730960, 64'd187209104, - 64'd30017622016, - 64'd15389016064, - 64'd408988352, 64'd173341968, - 64'd22354171904, - 64'd15248207872, - 64'd550607616, 64'd158774256, - 64'd14785753088, - 64'd15009643520, - 64'd683892544, 64'd143625904, - 64'd7360073728, - 64'd14678099968, - 64'd808224960, 64'd128016848, - 64'd122326760, - 64'd14258824192, - 64'd923066752, 64'd112066168, 64'd6885020160, - 64'd13757478912, - 64'd1027960576, 64'd95891384, 64'd13622423552, - 64'd13180087296, - 64'd1122530432, 64'd79607672, 64'd20053434368, - 64'd12532989952, - 64'd1206481152, 64'd63327192, 64'd26144839680, - 64'd11822783488, - 64'd1279598592, 64'd47158456, 64'd31866779648, - 64'd11056274432, - 64'd1341747456, 64'd31205682, 64'd37192835072, - 64'd10240421888, - 64'd1392870272, 64'd15568271, 64'd42100101120, - 64'd9382290432, - 64'd1432985088, 64'd340284, 64'd46569213952, - 64'd8488998400, - 64'd1462182656, - 64'd14390004, 64'd50584375296, - 64'd7567664640, - 64'd1480623872, - 64'd28540510, 64'd54133334016, - 64'd6625367552, - 64'd1488536064, - 64'd42035688, 64'd57207365632, - 64'd5669093376, - 64'd1486209792, - 64'd54806824, 64'd59801194496, - 64'd4705696256, - 64'd1473994240, - 64'd66792264, 64'd61912944640, - 64'd3741853952, - 64'd1452293376, - 64'd77937600, 64'd63544012800, - 64'd2784031744, - 64'd1421561344, - 64'd88195824, 64'd64698974208, - 64'd1838443904, - 64'd1382297856, - 64'd97527336, 64'd65385447424, - 64'd911020864, - 64'd1335043584, - 64'd105900048, 64'd65613926400, - 64'd7379710, - 64'd1280374656, - 64'd113289296, 64'd65397641216, 64'd867204224, - 64'd1218898048, - 64'd119677792, 64'd64752361472, 64'd1707821056, - 64'd1151246848, - 64'd125055480, 64'd63696216064, 64'd2509947136, - 64'd1078074240, - 64'd129419384, 64'd62249496576, 64'd3269463296, - 64'd1000049600, - 64'd132773400, 64'd60434452480, 64'd3982668544, - 64'd917852672, - 64'd135128032, 64'd58275078144, 64'd4646291968, - 64'd832168896, - 64'd136500128, 64'd55796891648, 64'd5257499648, - 64'd743684992, - 64'd136912544, 64'd53026709504, 64'd5813900800, - 64'd653083904, - 64'd136393792, 64'd49992445952, 64'd6313548288, - 64'd561040576, - 64'd134977664, 64'd46722871296, 64'd6754936320, - 64'd468217632, - 64'd132702888, 64'd43247403008, 64'd7136999424, - 64'd375261408, - 64'd129612640, 64'd39595872256, 64'd7459101696, - 64'd282798048, - 64'd125754136, 64'd35798339584, 64'd7721029120, - 64'd191430208, - 64'd121178200, 64'd31884855296, 64'd7922977280, - 64'd101733480, - 64'd115938792, 64'd27885277184, 64'd8065535488, - 64'd14253701, - 64'd110092552, 64'd23829073920, 64'd8149671936, 64'd70495888, - 64'd103698320, 64'd19745140736, 64'd8176712704, 64'd152036944, - 64'd96816696, 64'd15661621248, 64'd8148323328, 64'd229928128, - 64'd89509568, 64'd11605748736, 64'd8066485760, 64'd303766784, - 64'd81839656, 64'd7603688960, 64'd7933474816, 64'd373190432, - 64'd73870048, 64'd3680404224, 64'd7751833600, 64'd437877920, - 64'd65663800, - 64'd140476864, 64'd7524347392, 64'd497550080, - 64'd57283504, - 64'd3836774656, 64'd7254018048, 64'd551970432, - 64'd48790868, - 64'd7387857920, 64'd6944036352, 64'd600945152, - 64'd40246348, - 64'd10774731776, 64'd6597754880, 64'd644323200, - 64'd31708794, - 64'd13980114944, 64'd6218660352, 64'd681995840, - 64'd23235080, - 64'd16988492800, 64'd5810344448, 64'd713896000, - 64'd14879819, - 64'd19786172416, 64'd5376479744, 64'd739997248, - 64'd6695052, - 64'd22361307136, 64'd4920788992, 64'd760312896, 64'd1270005, - 64'd24703920128, 64'd4447020544, 64'd774894464, 64'd8969208, - 64'd26805911552, 64'd3958922496, 64'd783830144, 64'd16359686, - 64'd28661049344, 64'd3460217344, 64'd787242880, 64'd23402022, - 64'd30264948736, 64'd2954577408, 64'd785288704, 64'd30060408, - 64'd31615045632, 64'd2445602560, 64'd778154368, 64'd36302760, - 64'd32710555648, 64'd1936798720, 64'd766055168, 64'd42100824, - 64'd33552416768, 64'd1431556480, 64'd749232704, 64'd47430228, - 64'd34143229952, 64'd933133504, 64'd727952128, 64'd52270520, - 64'd34487185408, 64'd444635872, 64'd702499968, 64'd56605188, - 64'd34589990912, - 64'd30996946, 64'd673181248, 64'd60421624, - 64'd34458779648, - 64'd491006656, 64'd640316992, 64'd63711108, - 64'd34102003712, - 64'd932828672, 64'd604241408, 64'd66468712, - 64'd33529362432, - 64'd1354102784, 64'd565299456, 64'd68693224, - 64'd32751673344, - 64'd1752682880, 64'd523844032, 64'd70387048, - 64'd31780775936, - 64'd2126643328, 64'd480233312, 64'd71556032, - 64'd30629410816, - 64'd2474285568, 64'd434828384, 64'd72209368, - 64'd29311117312, - 64'd2794141952, 64'd387990528, 64'd72359368, - 64'd27840104448, - 64'd3084977920, 64'd340078944, 64'd72021344, - 64'd26231142400, - 64'd3345792256, 64'd291448352, 64'd71213336, - 64'd24499443712, - 64'd3575817216, 64'd242446768, 64'd69955968, - 64'd22660548608, - 64'd3774514944, 64'd193413440, 64'd68272184, - 64'd20730206208, - 64'd3941574912, 64'd144676800, 64'd66187028, - 64'd18724265984, - 64'd4076907264, 64'd96552704, 64'd63727432, - 64'd16658572288, - 64'd4180636928, 64'd49342632, 64'd60921944, - 64'd14548849664, - 64'd4253096448, 64'd3332228, 64'd57800504, - 64'd12410608640, - 64'd4294816000, - 64'd41210148, 64'd54394188, - 64'd10259047424, - 64'd4306513408, - 64'd84034640, 64'd50734972, - 64'd8108961280, - 64'd4289084160, - 64'd124910944, 64'd46855484, - 64'd5974653440, - 64'd4243589120, - 64'd163629248, 64'd42788764};


endpackage
`endif

