`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam N = 4;
	localparam M = 4;
	localparam real Lfr[0:3] = {0.98591065, 0.98591065, 0.9699685, 0.9699685};
	localparam real Lfi[0:3] = {0.059811182, -0.059811182, 0.023870276, -0.023870276};
	localparam real Lbr[0:3] = {0.98591065, 0.98591065, 0.9699685, 0.9699685};
	localparam real Lbi[0:3] = {0.059811182, -0.059811182, 0.023870276, -0.023870276};
	localparam real Wfr[0:3] = {-3.2207987e-05, -3.2207987e-05, 9.544637e-06, 9.544637e-06};
	localparam real Wfi[0:3] = {-1.418066e-06, 1.418066e-06, 1.8536752e-05, -1.8536752e-05};
	localparam real Wbr[0:3] = {3.2207987e-05, 3.2207987e-05, -9.544637e-06, -9.544637e-06};
	localparam real Wbi[0:3] = {1.418066e-06, -1.418066e-06, -1.8536752e-05, 1.8536752e-05};
	localparam real Ffr[0:3][0:79] = '{
		'{-94.38814, -11.340327, 1.5996957, -0.021420214, -99.80632, -10.3296995, 1.6094346, -0.02980436, -104.71543, -9.30473, 1.6128588, -0.037871376, -109.10935, -8.269639, 1.6101094, -0.045598533, -112.98406, -7.2285824, 1.6013476, -0.052964948, -116.33761, -6.1856356, 1.5867531, -0.05995162, -119.17004, -5.1447835, 1.5665233, -0.06654142, -121.483376, -4.1099052, 1.5408722, -0.072719164, -123.281555, -3.0847619, 1.5100288, -0.07847157, -124.57036, -2.0729873, 1.4742365, -0.08378731, -125.357346, -1.0780754, 1.433751, -0.08865695, -125.651794, -0.103371456, 1.3888398, -0.093073, -125.46461, 0.84793735, 1.3397804, -0.09702986, -124.80825, 1.7728299, 1.2868594, -0.10052378, -123.69665, 2.6684585, 1.2303708, -0.10355287, -122.14511, 3.5321555, 1.1706148, -0.10611705, -120.17023, 4.3614388, 1.107897, -0.10821796, -117.78979, 5.154017, 1.0425265, -0.10985899, -115.022675, 5.907793, 0.9748146, -0.11104516, -111.88877, 6.620868, 0.9050743, -0.11178308},
		'{-94.38814, -11.340327, 1.5996957, -0.021420214, -99.80632, -10.3296995, 1.6094346, -0.02980436, -104.71543, -9.30473, 1.6128588, -0.037871376, -109.10935, -8.269639, 1.6101094, -0.045598533, -112.98406, -7.2285824, 1.6013476, -0.052964948, -116.33761, -6.1856356, 1.5867531, -0.05995162, -119.17004, -5.1447835, 1.5665233, -0.06654142, -121.483376, -4.1099052, 1.5408722, -0.072719164, -123.281555, -3.0847619, 1.5100288, -0.07847157, -124.57036, -2.0729873, 1.4742365, -0.08378731, -125.357346, -1.0780754, 1.433751, -0.08865695, -125.651794, -0.103371456, 1.3888398, -0.093073, -125.46461, 0.84793735, 1.3397804, -0.09702986, -124.80825, 1.7728299, 1.2868594, -0.10052378, -123.69665, 2.6684585, 1.2303708, -0.10355287, -122.14511, 3.5321555, 1.1706148, -0.10611705, -120.17023, 4.3614388, 1.107897, -0.10821796, -117.78979, 5.154017, 1.0425265, -0.10985899, -115.022675, 5.907793, 0.9748146, -0.11104516, -111.88877, 6.620868, 0.9050743, -0.11178308},
		'{93.38552, 11.229796, -1.5223757, 0.26254022, 98.76348, 10.2888155, -1.4183407, 0.25036135, 103.680984, 9.387826, -1.3183138, 0.2385276, 108.15778, 8.525811, -1.2222077, 0.22703615, 112.21311, 7.7017555, -1.1299337, 0.21588388, 115.865685, 6.914648, -1.0414033, 0.20506734, 119.13373, 6.1634817, -0.9565275, 0.19458275, 122.03497, 5.447257, -0.87521684, 0.1844261, 124.58663, 4.76498, -0.79738235, 0.17459312, 126.80543, 4.115666, -0.7229347, 0.16507934, 128.70761, 3.498339, -0.6517852, 0.15588003, 130.30893, 2.9120338, -0.58384514, 0.14699031, 131.62463, 2.3557954, -0.5190266, 0.13840513, 132.66956, 1.8286806, -0.45724198, 0.13011928, 133.45801, 1.3297591, -0.39840454, 0.12212742, 134.00385, 0.858113, -0.3424281, 0.11442408, 134.3205, 0.4128385, -0.28922746, 0.10700369, 134.42091, -0.0069543985, -0.23871827, 0.09986059, 134.31763, -0.40214083, -0.19081716, 0.092989065, 134.02272, -0.7735809, -0.14544182, 0.08638329},
		'{93.38552, 11.229796, -1.5223757, 0.26254022, 98.76348, 10.2888155, -1.4183407, 0.25036135, 103.680984, 9.387826, -1.3183138, 0.2385276, 108.15778, 8.525811, -1.2222077, 0.22703615, 112.21311, 7.7017555, -1.1299337, 0.21588388, 115.865685, 6.914648, -1.0414033, 0.20506734, 119.13373, 6.1634817, -0.9565275, 0.19458275, 122.03497, 5.447257, -0.87521684, 0.1844261, 124.58663, 4.76498, -0.79738235, 0.17459312, 126.80543, 4.115666, -0.7229347, 0.16507934, 128.70761, 3.498339, -0.6517852, 0.15588003, 130.30893, 2.9120338, -0.58384514, 0.14699031, 131.62463, 2.3557954, -0.5190266, 0.13840513, 132.66956, 1.8286806, -0.45724198, 0.13011928, 133.45801, 1.3297591, -0.39840454, 0.12212742, 134.00385, 0.858113, -0.3424281, 0.11442408, 134.3205, 0.4128385, -0.28922746, 0.10700369, 134.42091, -0.0069543985, -0.23871827, 0.09986059, 134.31763, -0.40214083, -0.19081716, 0.092989065, 134.02272, -0.7735809, -0.14544182, 0.08638329}};
	localparam real Ffi[0:3][0:79] = '{
		'{112.82257, -14.225602, -0.53965706, 0.14522274, 105.58751, -14.703451, -0.43637398, 0.14189547, 98.13032, -15.114121, -0.33396357, 0.13811363, 90.48457, -15.457701, -0.23279127, 0.13390256, 82.68375, -15.734529, -0.13320884, 0.12928867, 74.76108, -15.945189, -0.035553526, 0.12429918, 66.74946, -16.090504, 0.05985298, 0.11896212, 58.6813, -16.171515, 0.15270531, 0.1133061, 50.58846, -16.189487, 0.24271518, 0.10736027, 42.502083, -16.145891, 0.3296121, 0.10115416, 34.452557, -16.042395, 0.4131439, 0.09471755, 26.469374, -15.880849, 0.49307734, 0.08808037, 18.581055, -15.663281, 0.56919837, 0.081272565, 10.815074, -15.39188, 0.6413126, 0.07432402, 3.197768, -15.068984, 0.7092455, 0.0672644, -4.2457294, -14.697068, 0.77284265, 0.06012307, -11.491553, -14.278734, 0.8319697, 0.05292899, -18.517168, -13.816693, 0.8865124, 0.045710612, -25.30142, -13.313758, 0.9363768, 0.038495783, -31.824583, -12.772824, 0.9814887, 0.03131166},
		'{-112.82257, 14.225602, 0.53965706, -0.14522274, -105.58751, 14.703451, 0.43637398, -0.14189547, -98.13032, 15.114121, 0.33396357, -0.13811363, -90.48457, 15.457701, 0.23279127, -0.13390256, -82.68375, 15.734529, 0.13320884, -0.12928867, -74.76108, 15.945189, 0.035553526, -0.12429918, -66.74946, 16.090504, -0.05985298, -0.11896212, -58.6813, 16.171515, -0.15270531, -0.1133061, -50.58846, 16.189487, -0.24271518, -0.10736027, -42.502083, 16.145891, -0.3296121, -0.10115416, -34.452557, 16.042395, -0.4131439, -0.09471755, -26.469374, 15.880849, -0.49307734, -0.08808037, -18.581055, 15.663281, -0.56919837, -0.081272565, -10.815074, 15.39188, -0.6413126, -0.07432402, -3.197768, 15.068984, -0.7092455, -0.0672644, 4.2457294, 14.697068, -0.77284265, -0.06012307, 11.491553, 14.278734, -0.8319697, -0.05292899, 18.517168, 13.816693, -0.8865124, -0.045710612, 25.30142, 13.313758, -0.9363768, -0.038495783, 31.824583, 12.772824, -0.9814887, -0.03131166},
		'{-342.78888, 25.292248, -2.443028, 0.17990588, -330.26526, 24.800743, -2.4059997, 0.18076995, -317.98938, 24.301537, -2.3676, 0.18131734, -305.9648, 23.795815, -2.327966, 0.18156584, -294.19446, 23.284702, -2.287228, 0.18153255, -282.6808, 22.769272, -2.245511, 0.18123406, -271.42572, 22.25053, -2.2029335, 0.18068634, -260.43063, 21.729437, -2.1596086, 0.1799048, -249.6965, 21.206898, -2.115644, 0.1789043, -239.22383, 20.683764, -2.0711417, 0.17769912, -229.0127, 20.160841, -2.0261989, 0.17630303, -219.0628, 19.638887, -1.9809074, 0.17472929, -209.3735, 19.118612, -1.9353544, 0.1729906, -199.94379, 18.600685, -1.889622, 0.1710992, -190.77232, 18.08573, -1.8437883, 0.16906682, -181.85745, 17.57433, -1.7979265, 0.1669047, -173.1973, 17.06703, -1.752106, 0.16462363, -164.78966, 16.564335, -1.7063916, 0.16223395, -156.63211, 16.066717, -1.6608443, 0.15974551, -148.72202, 15.57461, -1.6155214, 0.15716779},
		'{342.78888, -25.292248, 2.443028, -0.17990588, 330.26526, -24.800743, 2.4059997, -0.18076995, 317.98938, -24.301537, 2.3676, -0.18131734, 305.9648, -23.795815, 2.327966, -0.18156584, 294.19446, -23.284702, 2.287228, -0.18153255, 282.6808, -22.769272, 2.245511, -0.18123406, 271.42572, -22.25053, 2.2029335, -0.18068634, 260.43063, -21.729437, 2.1596086, -0.1799048, 249.6965, -21.206898, 2.115644, -0.1789043, 239.22383, -20.683764, 2.0711417, -0.17769912, 229.0127, -20.160841, 2.0261989, -0.17630303, 219.0628, -19.638887, 1.9809074, -0.17472929, 209.3735, -19.118612, 1.9353544, -0.1729906, 199.94379, -18.600685, 1.889622, -0.1710992, 190.77232, -18.08573, 1.8437883, -0.16906682, 181.85745, -17.57433, 1.7979265, -0.1669047, 173.1973, -17.06703, 1.752106, -0.16462363, 164.78966, -16.564335, 1.7063916, -0.16223395, 156.63211, -16.066717, 1.6608443, -0.15974551, 148.72202, -15.57461, 1.6155214, -0.15716779}};
	localparam real Fbr[0:3][0:79] = '{
		'{94.38814, -11.340327, -1.5996957, -0.021420214, 99.80632, -10.3296995, -1.6094346, -0.02980436, 104.71543, -9.30473, -1.6128588, -0.037871376, 109.10935, -8.269639, -1.6101094, -0.045598533, 112.98406, -7.2285824, -1.6013476, -0.052964948, 116.33761, -6.1856356, -1.5867531, -0.05995162, 119.17004, -5.1447835, -1.5665233, -0.06654142, 121.483376, -4.1099052, -1.5408722, -0.072719164, 123.281555, -3.0847619, -1.5100288, -0.07847157, 124.57036, -2.0729873, -1.4742365, -0.08378731, 125.357346, -1.0780754, -1.433751, -0.08865695, 125.651794, -0.103371456, -1.3888398, -0.093073, 125.46461, 0.84793735, -1.3397804, -0.09702986, 124.80825, 1.7728299, -1.2868594, -0.10052378, 123.69665, 2.6684585, -1.2303708, -0.10355287, 122.14511, 3.5321555, -1.1706148, -0.10611705, 120.17023, 4.3614388, -1.107897, -0.10821796, 117.78979, 5.154017, -1.0425265, -0.10985899, 115.022675, 5.907793, -0.9748146, -0.11104516, 111.88877, 6.620868, -0.9050743, -0.11178308},
		'{94.38814, -11.340327, -1.5996957, -0.021420214, 99.80632, -10.3296995, -1.6094346, -0.02980436, 104.71543, -9.30473, -1.6128588, -0.037871376, 109.10935, -8.269639, -1.6101094, -0.045598533, 112.98406, -7.2285824, -1.6013476, -0.052964948, 116.33761, -6.1856356, -1.5867531, -0.05995162, 119.17004, -5.1447835, -1.5665233, -0.06654142, 121.483376, -4.1099052, -1.5408722, -0.072719164, 123.281555, -3.0847619, -1.5100288, -0.07847157, 124.57036, -2.0729873, -1.4742365, -0.08378731, 125.357346, -1.0780754, -1.433751, -0.08865695, 125.651794, -0.103371456, -1.3888398, -0.093073, 125.46461, 0.84793735, -1.3397804, -0.09702986, 124.80825, 1.7728299, -1.2868594, -0.10052378, 123.69665, 2.6684585, -1.2303708, -0.10355287, 122.14511, 3.5321555, -1.1706148, -0.10611705, 120.17023, 4.3614388, -1.107897, -0.10821796, 117.78979, 5.154017, -1.0425265, -0.10985899, 115.022675, 5.907793, -0.9748146, -0.11104516, 111.88877, 6.620868, -0.9050743, -0.11178308},
		'{-93.38552, 11.229796, 1.5223757, 0.26254022, -98.76348, 10.2888155, 1.4183407, 0.25036135, -103.680984, 9.387826, 1.3183138, 0.2385276, -108.15778, 8.525811, 1.2222077, 0.22703615, -112.21311, 7.7017555, 1.1299337, 0.21588388, -115.865685, 6.914648, 1.0414033, 0.20506734, -119.13373, 6.1634817, 0.9565275, 0.19458275, -122.03497, 5.447257, 0.87521684, 0.1844261, -124.58663, 4.76498, 0.79738235, 0.17459312, -126.80543, 4.115666, 0.7229347, 0.16507934, -128.70761, 3.498339, 0.6517852, 0.15588003, -130.30893, 2.9120338, 0.58384514, 0.14699031, -131.62463, 2.3557954, 0.5190266, 0.13840513, -132.66956, 1.8286806, 0.45724198, 0.13011928, -133.45801, 1.3297591, 0.39840454, 0.12212742, -134.00385, 0.858113, 0.3424281, 0.11442408, -134.3205, 0.4128385, 0.28922746, 0.10700369, -134.42091, -0.0069543985, 0.23871827, 0.09986059, -134.31763, -0.40214083, 0.19081716, 0.092989065, -134.02272, -0.7735809, 0.14544182, 0.08638329},
		'{-93.38552, 11.229796, 1.5223757, 0.26254022, -98.76348, 10.2888155, 1.4183407, 0.25036135, -103.680984, 9.387826, 1.3183138, 0.2385276, -108.15778, 8.525811, 1.2222077, 0.22703615, -112.21311, 7.7017555, 1.1299337, 0.21588388, -115.865685, 6.914648, 1.0414033, 0.20506734, -119.13373, 6.1634817, 0.9565275, 0.19458275, -122.03497, 5.447257, 0.87521684, 0.1844261, -124.58663, 4.76498, 0.79738235, 0.17459312, -126.80543, 4.115666, 0.7229347, 0.16507934, -128.70761, 3.498339, 0.6517852, 0.15588003, -130.30893, 2.9120338, 0.58384514, 0.14699031, -131.62463, 2.3557954, 0.5190266, 0.13840513, -132.66956, 1.8286806, 0.45724198, 0.13011928, -133.45801, 1.3297591, 0.39840454, 0.12212742, -134.00385, 0.858113, 0.3424281, 0.11442408, -134.3205, 0.4128385, 0.28922746, 0.10700369, -134.42091, -0.0069543985, 0.23871827, 0.09986059, -134.31763, -0.40214083, 0.19081716, 0.092989065, -134.02272, -0.7735809, 0.14544182, 0.08638329}};
	localparam real Fbi[0:3][0:79] = '{
		'{-112.82257, -14.225602, 0.53965706, 0.14522274, -105.58751, -14.703451, 0.43637398, 0.14189547, -98.13032, -15.114121, 0.33396357, 0.13811363, -90.48457, -15.457701, 0.23279127, 0.13390256, -82.68375, -15.734529, 0.13320884, 0.12928867, -74.76108, -15.945189, 0.035553526, 0.12429918, -66.74946, -16.090504, -0.05985298, 0.11896212, -58.6813, -16.171515, -0.15270531, 0.1133061, -50.58846, -16.189487, -0.24271518, 0.10736027, -42.502083, -16.145891, -0.3296121, 0.10115416, -34.452557, -16.042395, -0.4131439, 0.09471755, -26.469374, -15.880849, -0.49307734, 0.08808037, -18.581055, -15.663281, -0.56919837, 0.081272565, -10.815074, -15.39188, -0.6413126, 0.07432402, -3.197768, -15.068984, -0.7092455, 0.0672644, 4.2457294, -14.697068, -0.77284265, 0.06012307, 11.491553, -14.278734, -0.8319697, 0.05292899, 18.517168, -13.816693, -0.8865124, 0.045710612, 25.30142, -13.313758, -0.9363768, 0.038495783, 31.824583, -12.772824, -0.9814887, 0.03131166},
		'{112.82257, 14.225602, -0.53965706, -0.14522274, 105.58751, 14.703451, -0.43637398, -0.14189547, 98.13032, 15.114121, -0.33396357, -0.13811363, 90.48457, 15.457701, -0.23279127, -0.13390256, 82.68375, 15.734529, -0.13320884, -0.12928867, 74.76108, 15.945189, -0.035553526, -0.12429918, 66.74946, 16.090504, 0.05985298, -0.11896212, 58.6813, 16.171515, 0.15270531, -0.1133061, 50.58846, 16.189487, 0.24271518, -0.10736027, 42.502083, 16.145891, 0.3296121, -0.10115416, 34.452557, 16.042395, 0.4131439, -0.09471755, 26.469374, 15.880849, 0.49307734, -0.08808037, 18.581055, 15.663281, 0.56919837, -0.081272565, 10.815074, 15.39188, 0.6413126, -0.07432402, 3.197768, 15.068984, 0.7092455, -0.0672644, -4.2457294, 14.697068, 0.77284265, -0.06012307, -11.491553, 14.278734, 0.8319697, -0.05292899, -18.517168, 13.816693, 0.8865124, -0.045710612, -25.30142, 13.313758, 0.9363768, -0.038495783, -31.824583, 12.772824, 0.9814887, -0.03131166},
		'{342.78888, 25.292248, 2.443028, 0.17990588, 330.26526, 24.800743, 2.4059997, 0.18076995, 317.98938, 24.301537, 2.3676, 0.18131734, 305.9648, 23.795815, 2.327966, 0.18156584, 294.19446, 23.284702, 2.287228, 0.18153255, 282.6808, 22.769272, 2.245511, 0.18123406, 271.42572, 22.25053, 2.2029335, 0.18068634, 260.43063, 21.729437, 2.1596086, 0.1799048, 249.6965, 21.206898, 2.115644, 0.1789043, 239.22383, 20.683764, 2.0711417, 0.17769912, 229.0127, 20.160841, 2.0261989, 0.17630303, 219.0628, 19.638887, 1.9809074, 0.17472929, 209.3735, 19.118612, 1.9353544, 0.1729906, 199.94379, 18.600685, 1.889622, 0.1710992, 190.77232, 18.08573, 1.8437883, 0.16906682, 181.85745, 17.57433, 1.7979265, 0.1669047, 173.1973, 17.06703, 1.752106, 0.16462363, 164.78966, 16.564335, 1.7063916, 0.16223395, 156.63211, 16.066717, 1.6608443, 0.15974551, 148.72202, 15.57461, 1.6155214, 0.15716779},
		'{-342.78888, -25.292248, -2.443028, -0.17990588, -330.26526, -24.800743, -2.4059997, -0.18076995, -317.98938, -24.301537, -2.3676, -0.18131734, -305.9648, -23.795815, -2.327966, -0.18156584, -294.19446, -23.284702, -2.287228, -0.18153255, -282.6808, -22.769272, -2.245511, -0.18123406, -271.42572, -22.25053, -2.2029335, -0.18068634, -260.43063, -21.729437, -2.1596086, -0.1799048, -249.6965, -21.206898, -2.115644, -0.1789043, -239.22383, -20.683764, -2.0711417, -0.17769912, -229.0127, -20.160841, -2.0261989, -0.17630303, -219.0628, -19.638887, -1.9809074, -0.17472929, -209.3735, -19.118612, -1.9353544, -0.1729906, -199.94379, -18.600685, -1.889622, -0.1710992, -190.77232, -18.08573, -1.8437883, -0.16906682, -181.85745, -17.57433, -1.7979265, -0.1669047, -173.1973, -17.06703, -1.752106, -0.16462363, -164.78966, -16.564335, -1.7063916, -0.16223395, -156.63211, -16.066717, -1.6608443, -0.15974551, -148.72202, -15.57461, -1.6155214, -0.15716779}};
	localparam real hf[0:1199] = {0.02089113, -3.3151082e-05, -4.3065935e-05, 1.3363545e-07, 0.020857995, -9.934768e-05, -4.2787167e-05, 3.9975208e-07, 0.020791832, -0.00016522867, -4.223146e-05, 6.624789e-07, 0.020692853, -0.00023058585, -4.1402196e-05, 9.197127e-07, 0.020561367, -0.00029521363, -4.030422e-05, 1.1694873e-06, 0.020397792, -0.00035890998, -3.8943755e-05, 1.4099754e-06, 0.020202644, -0.00042147728, -3.7328326e-05, 1.63949e-06, 0.019976534, -0.0004827232, -3.5466684e-05, 1.8564855e-06, 0.01972017, -0.0005424616, -3.336872e-05, 2.0595573e-06, 0.019434351, -0.0006005129, -3.1045372e-05, 2.247443e-06, 0.019119965, -0.00065670535, -2.850855e-05, 2.4190206e-06, 0.018777981, -0.00071087515, -2.5771038e-05, 2.573307e-06, 0.018409451, -0.0007628674, -2.2846416e-05, 2.7094582e-06, 0.0180155, -0.00081253634, -1.9748964e-05, 2.8267657e-06, 0.017597325, -0.0008597462, -1.649358e-05, 2.9246546e-06, 0.017156184, -0.00090437126, -1.309568e-05, 3.0026804e-06, 0.016693402, -0.0009462965, -9.5711275e-06, 3.0605268e-06, 0.016210355, -0.0009854177, -5.936136e-06, 3.0980007e-06, 0.015708467, -0.0010216419, -2.2071874e-06, 3.1150287e-06, 0.015189208, -0.0010548875, 1.5990514e-06, 3.1116538e-06, 0.014654087, -0.0010850846, 5.465811e-06, 3.0880294e-06, 0.014104641, -0.0011121746, 9.376297e-06, 3.0444157e-06, 0.013542437, -0.001136111, 1.3313769e-05, 2.9811733e-06, 0.012969061, -0.0011568589, 1.7261615e-05, 2.89876e-06, 0.012386113, -0.0011743947, 2.1203417e-05, 2.7977223e-06, 0.011795203, -0.0011887072, 2.5123034e-05, 2.6786931e-06, 0.011197943, -0.0011997957, 2.9004652e-05, 2.5423833e-06, 0.010595943, -0.0012076716, 3.2832853e-05, 2.3895775e-06, 0.009990803, -0.0012123566, 3.659268e-05, 2.221127e-06, 0.009384112, -0.0012138837, 4.0269675e-05, 2.0379443e-06, 0.008777439, -0.0012122962, 4.3849952e-05, 1.8409968e-06, 0.008172326, -0.0012076475, 4.732023e-05, 1.6313006e-06, 0.0075702905, -0.0012000008, 5.0667884e-05, 1.4099147e-06, 0.006972813, -0.0011894285, 5.3880976e-05, 1.1779345e-06, 0.006381336, -0.0011760121, 5.6948305e-05, 9.364856e-07, 0.00579726, -0.0011598415, 5.9859427e-05, 6.867187e-07, 0.0052219373, -0.0011410147, 6.260469e-05, 4.2980258e-07, 0.0046566706, -0.0011196368, 6.5175256e-05, 1.6691912e-07, 0.0041027074, -0.0010958203, 6.7563116e-05, -1.00742795e-07, 0.0035612374, -0.0010696838, 6.976111e-05, -3.7199266e-07, 0.0030333898, -0.0010413518, 7.176296e-05, -6.456437e-07, 0.0025202301, -0.0010109541, 7.356322e-05, -9.2051806e-07, 0.002022758, -0.0009786253, 7.515736e-05, -1.1954519e-06, 0.0015419039, -0.000944504, 7.65417e-05, -1.4693001e-06, 0.0010785293, -0.0009087323, 7.7713434e-05, -1.7409408e-06, 0.00063342287, -0.00087145536, 7.867064e-05, -2.0092798e-06, 0.00020730059, -0.00083282066, 7.941223e-05, -2.273255e-06, -0.000199196, -0.0007929776, 7.993798e-05, -2.531839e-06, -0.0005855002, -0.0007520764, 8.024848e-05, -2.7840447e-06, -0.00095112086, -0.00071026833, 8.034514e-05, -3.028927e-06, -0.0012956422, -0.0006677045, 8.023015e-05, -3.2655869e-06, -0.0016187241, -0.0006245356, 7.990647e-05, -3.493173e-06, -0.0019201015, -0.00058091135, 7.937779e-05, -3.7108857e-06, -0.002199584, -0.0005369799, 7.86485e-05, -3.9179786e-06, -0.002457054, -0.00049288716, 7.772369e-05, -4.1137596e-06, -0.0026924678, -0.00044877693, 7.660907e-05, -4.297595e-06, -0.0029058512, -0.00040478964, 7.5310956e-05, -4.4689077e-06, -0.0030973004, -0.0003610625, 7.383625e-05, -4.6271816e-06, -0.003266979, -0.00031772873, 7.219238e-05, -4.77196e-06, -0.0034151159, -0.00027491737, 7.038726e-05, -4.9028476e-06, -0.0035420037, -0.0002327528, 6.842926e-05, -5.01951e-06, -0.003647996, -0.00019135444, 6.632717e-05, -5.1216743e-06, -0.0037335046, -0.00015083635, 6.409014e-05, -5.209129e-06, -0.003798997, -0.00011130705, 6.172764e-05, -5.281723e-06, -0.0038449934, -7.286914e-05, 5.924944e-05, -5.3393655e-06, -0.003872064, -3.561914e-05, 5.666554e-05, -5.3820245e-06, -0.0038808254, 3.5276486e-07, 5.398614e-05, -5.4097272e-06, -0.003871938, 3.49629e-05, 5.12216e-05, -5.4225566e-06, -0.003846102, 6.813426e-05, 4.8382382e-05, -5.420651e-06, -0.003804055, 9.979662e-05, 4.547903e-05, -5.404204e-06, -0.0037465673, 0.00012988667, 4.2522115e-05, -5.373458e-06, -0.0036744396, 0.00015834805, 3.9522194e-05, -5.3287076e-06, -0.0035884988, 0.00018513142, 3.6489775e-05, -5.270295e-06, -0.003489595, 0.00021019446, 3.343528e-05, -5.198606e-06, -0.003378597, 0.0002335019, 3.0369003e-05, -5.1140705e-06, -0.0032563903, 0.0002550254, 2.7301081e-05, -5.017158e-06, -0.0031238724, 0.00027474365, 2.4241448e-05, -4.908377e-06, -0.00298195, 0.0002926421, 2.1199816e-05, -4.7882686e-06, -0.002831535, 0.00030871294, 1.8185634e-05, -4.657408e-06, -0.002673542, 0.000322955, 1.5208058e-05, -4.5163997e-06, -0.002508884, 0.0003353736, 1.2275935e-05, -4.365872e-06, -0.0023384704, 0.00034598025, 9.39776e-06, -4.2064794e-06, -0.002163203, 0.00035479266, 6.5816644e-06, -4.0388954e-06, -0.001983973, 0.0003618344, 3.83539e-06, -3.863811e-06, -0.0018016589, 0.00036713466, 1.1662675e-06, -3.6819313e-06, -0.0016171229, 0.00037072808, -1.4188005e-06, -3.4939735e-06, -0.0014312087, 0.00037265453, -3.9133556e-06, -3.3006627e-06, -0.0012447389, 0.0003729587, -6.3113976e-06, -3.1027296e-06, -0.0010585124, 0.00037168985, -8.607398e-06, -2.900908e-06, -0.00087330246, 0.00036890176, -1.0796308e-05, -2.6959303e-06, -0.00068985444, 0.00036465205, -1.2873567e-05, -2.4885273e-06, -0.00050888397, 0.00035900212, -1.4835111e-05, -2.2794236e-06, -0.00033107505, 0.00035201685, -1.6677372e-05, -2.0693353e-06, -0.00015707855, 0.00034376408, -1.8397284e-05, -1.8589683e-06, 1.2489361e-05, 0.00033431454, -1.9992282e-05, -1.6490147e-06, 0.0001770485, 0.00032374132, -2.1460299e-05, -1.4401517e-06, 0.0003360557, 0.0003121196, -2.2799763e-05, -1.2330385e-06, 0.000489006, 0.00029952647, -2.4009592e-05, -1.0283145e-06, 0.0006354331, 0.0002860403, -2.508919e-05, -8.265978e-07, 0.00077491056, 0.0002717408, -2.6038428e-05, -6.2848255e-07, 0.00090705155, 0.00025670833, -2.6857646e-05, -4.3453778e-07, 0.00103151, 0.0002410238, -2.7547636e-05, -2.4530576e-07, 0.00114798, 0.00022476834, -2.8109625e-05, -6.130047e-08, 0.0012561965, 0.00020802299, -2.8545266e-05, 1.1699363e-07, 0.0013559345, 0.0001908683, -2.8856623e-05, 2.8912274e-07, 0.0014470097, 0.00017338422, -2.9046143e-05, 4.5466476e-07, 0.0015292768, 0.00015564967, -2.9116654e-05, 6.132301e-07, 0.0016026304, 0.00013774236, -2.9071338e-05, 7.6446247e-07, 0.001667003, 0.00011973852, -2.8913702e-05, 9.080394e-07, 0.0017223652, 0.00010171263, -2.864758e-05, 1.0436728e-06, 0.001768724, 8.37372e-05, -2.8277087e-05, 1.1711089e-06, 0.0018061224, 6.588259e-05, -2.7806615e-05, 1.290129e-06, 0.0018346378, 4.8216738e-05, -2.7240796e-05, 1.400549e-06, 0.0018543813, 3.080503e-05, -2.65845e-05, 1.5022194e-06, 0.0018654956, 1.3710084e-05, -2.5842783e-05, 1.5950253e-06, 0.001868154, -3.008397e-06, -2.502089e-05, 1.6788858e-06, 0.0018625592, -1.9293771e-05, -2.412422e-05, 1.7537535e-06, 0.0018489413, -3.5092595e-05, -2.3158298e-05, 1.8196142e-06, 0.001827556, -5.0354738e-05, -2.2128765e-05, 1.876486e-06, 0.0017986838, -6.503348e-05, -2.1041336e-05, 1.924418e-06, 0.001762627, -7.908561e-05, -1.99018e-05, 1.963491e-06, 0.0017197091, -9.2471484e-05, -1.8715973e-05, 1.9938143e-06, 0.0016702726, -0.000105155086, -1.74897e-05, 2.0155262e-06, 0.0016146766, -0.00011710408, -1.6228809e-05, 2.0287923e-06, 0.0015532956, -0.00012828982, -1.4939109e-05, 2.0338043e-06, 0.0014865181, -0.00013868736, -1.362636e-05, 2.0307787e-06, 0.0014147433, -0.00014827549, -1.2296254e-05, 2.0199554e-06, 0.0013383805, -0.00015703666, -1.0954395e-05, 2.0015964e-06, 0.0012578468, -0.000164957, -9.606287e-06, 1.975984e-06, 0.0011735654, -0.00017202628, -8.257306e-06, 1.9434199e-06, 0.0010859636, -0.00017823778, -6.912691e-06, 1.9042225e-06, 0.0009954711, -0.00018358832, -5.577525e-06, 1.8587268e-06, 0.00090251875, -0.00018807813, -4.2567203e-06, 1.8072818e-06, 0.00080753595, -0.0001917108, -2.955006e-06, 1.750249e-06, 0.00071094977, -0.00019449311, -1.676913e-06, 1.688001e-06, 0.000613183, -0.000196435, -4.2676385e-07, 1.6209199e-06, 0.0005146528, -0.00019754937, 7.913391e-07, 1.5493953e-06, 0.00041576906, -0.00019785204, 1.9735228e-06, 1.4738231e-06, 0.0003169331, -0.00019736159, 3.1161526e-06, 1.3946036e-06, 0.00021853628, -0.00019609914, 4.215839e-06, 1.3121403e-06, 0.000120958815, -0.00019408834, 5.2694445e-06, 1.2268376e-06, 2.4568484e-05, -0.00019135511, 6.27409e-06, 1.1391004e-06, -7.0280425e-05, -0.00018792751, 7.227157e-06, 1.0493314e-06, -0.00016324816, -0.00018383561, 8.1262915e-06, 9.579305e-07, -0.0002540105, -0.00017911129, 8.969408e-06, 8.6529326e-07, -0.00034225947, -0.00017378808, 9.754686e-06, 7.7180914e-07, -0.00042770442, -0.00016790099, 1.0480577e-05, 6.778606e-07, -0.0005100724, -0.00016148636, 1.1145795e-05, 5.838219e-07, -0.00058910897, -0.00015458165, 1.1749322e-05, 4.900576e-07, -0.00066457863, -0.0001472253, 1.22904e-05, 3.9692156e-07, -0.0007362654, -0.00013945656, 1.27685325e-05, 3.047562e-07, -0.00080397294, -0.00013131526, 1.3183473e-05, 2.138912e-07, -0.0008675251, -0.00012284175, 1.3535224e-05, 1.2464257e-07, -0.00092676596, -0.00011407665, 1.3824031e-05, 3.7312006e-08, -0.0009815599, -0.000105060666, 1.4050373e-05, -4.781396e-08, -0.0010317914, -9.583455e-05, 1.4214956e-05, -1.3046464e-07, -0.001077366, -8.643882e-05, 1.4318705e-05, -2.103858e-07, -0.0011182086, -7.691369e-05, 1.4362755e-05, -2.8734019e-07, -0.0011542646, -6.729886e-05, 1.43484385e-05, -3.6110802e-07, -0.0011854989, -5.7633446e-05, 1.427728e-05, -4.3148725e-07, -0.0012118958, -4.7955797e-05, 1.4150984e-05, -4.9829407e-07, -0.0012334588, -3.8303377e-05, 1.3971419e-05, -5.61363e-07, -0.0012502094, -2.8712651e-05, 1.3740616e-05, -6.205469e-07, -0.0012621875, -1.9218973e-05, 1.3460747e-05, -6.7571756e-07, -0.0012694502, -9.856461e-06, 1.31341185e-05, -7.2676505e-07, -0.0012720713, -6.579164e-07, 1.276316e-05, -7.735982e-07, -0.0012701406, 8.345278e-06, 1.2350408e-05, -8.1614405e-07, -0.0012637634, 1.7123242e-05, 1.1898494e-05, -8.543481e-07, -0.0012530595, 2.5647678e-05, 1.1410139e-05, -8.881737e-07, -0.0012381624, 3.389193e-05, 1.0888131e-05, -9.176018e-07, -0.0012192184, 4.1831066e-05, 1.03353195e-05, -9.4263083e-07, -0.0011963861, 4.9441896e-05, 9.7546e-06, -9.632757e-07, -0.0011698348, 5.6703062e-05, 9.148904e-06, -9.795682e-07, -0.0011397444, 6.3595035e-05, 8.521183e-06, -9.915556e-07, -0.0011063041, 7.010016e-05, 7.874404e-06, -9.993003e-07, -0.0010697114, 7.6202705e-05, 7.2115313e-06, -1.0028796e-06, -0.0010301708, 8.1888815e-05, 6.535516e-06, -1.0023847e-06, -0.0009878939, 8.7146575e-05, 5.849289e-06, -9.979202e-07, -0.00094309734, 9.1965965e-05, 5.1557467e-06, -9.89603e-07, -0.0008960024, 9.6338896e-05, 4.457742e-06, -9.775619e-07, -0.0008468339, 0.00010025915, 3.7580744e-06, -9.619366e-07, -0.00079581945, 0.00010372239, 3.0594817e-06, -9.428773e-07, -0.00074318814, 0.000106726126, 2.36463e-06, -9.205432e-07, -0.00068917003, 0.000109269655, 1.6761053e-06, -8.9510223e-07, -0.00063399505, 0.00011135404, 9.964059e-07, -8.6673e-07, -0.00057789206, 0.00011298208, 3.2793542e-07, -8.356088e-07, -0.0005210883, 0.000114158225, -3.2700433e-07, -8.0192706e-07, -0.00046380822, 0.000114888535, -9.662197e-07, -7.658782e-07, -0.00040627285, 0.000115180614, -1.5876305e-06, -7.2765994e-07, -0.00034869916, 0.00011504354, -2.1892758e-06, -6.8747323e-07, -0.00029129916, 0.000114487826, -2.7693175e-06, -6.455217e-07, -0.00023427921, 0.00011352528, -3.3260449e-06, -6.020107e-07, -0.00017783955, 0.000112169015, -3.8578783e-06, -5.571463e-07, -0.00012217351, 0.000110433284, -4.363371e-06, -5.111347e-07, -6.746702e-05, 0.00010833344, -4.841212e-06, -4.6418145e-07, -1.38980895e-05, 0.00010588588, -5.2902283e-06, -4.164905e-07, 3.8363713e-05, 0.00010310789, -5.7093844e-06, -3.682637e-07, 8.915767e-05, 0.00010001759, -6.097784e-06, -3.1969986e-07, 0.00013833233, 9.6633885e-05, -6.4546707e-06, -2.7099426e-07, 0.00018574584, 9.2976305e-05, -6.779425e-06, -2.2233787e-07, 0.00023126627, 8.906495e-05, -7.0715655e-06, -1.7391679e-07, 0.00027477185, 8.492043e-05, -7.330747e-06, -1.2591161e-07, 0.00031615124, 8.0563696e-05, -7.5567577e-06, -7.8496946e-08, 0.00035530367, 7.6016026e-05, -7.749518e-06, -3.1840855e-08, 0.00039213896, 7.129892e-05, -7.909074e-06, 1.38956295e-08, 0.00042657787, 6.643398e-05, -8.035602e-06, 5.855892e-08, 0.00045855186, 6.1442865e-05, -8.129394e-06, 1.020033e-07, 0.00048800325, 5.634719e-05, -8.190864e-06, 1.4409123e-07, 0.0005148851, 5.116844e-05, -8.220535e-06, 1.8469376e-07, 0.0005391613, 4.5927904e-05, -8.219043e-06, 2.236907e-07, 0.0005608062, 4.06466e-05, -8.187122e-06, 2.6097098e-07, 0.00057980453, 3.534518e-05, -8.125607e-06, 2.964327e-07, 0.00059615134, 3.00439e-05, -8.035425e-06, 3.299834e-07, 0.0006098517, 2.4762514e-05, -7.917587e-06, 3.6154026e-07, 0.0006209203, 1.9520232e-05, -7.773189e-06, 3.9102994e-07, 0.00062938145, 1.4335658e-05, -7.603398e-06, 4.183888e-07, 0.0006352685, 9.226734e-06, -7.4094505e-06, 4.4356287e-07, 0.00063862366, 4.210683e-06, -7.192644e-06, 4.6650783e-07, 0.0006394974, -6.9603163e-07, -6.954332e-06, 4.8718886e-07, 0.0006379484, -5.4777533e-06, -6.6959183e-06, 5.055807e-07, 0.0006340429, -1.0119673e-05, -6.4188466e-06, 5.216673e-07, 0.0006278543, -1.460786e-05, -6.1245987e-06, 5.3544187e-07, 0.0006194628, -1.89293e-05, -5.8146848e-06, 5.469065e-07, 0.0006089548, -2.3071916e-05, -5.490638e-06, 5.560721e-07, 0.0005964225, -2.7024593e-05, -5.1540096e-06, 5.62958e-07, 0.00058196357, -3.0777202e-05, -4.806359e-06, 5.6759166e-07, 0.0005656802, -3.43206e-05, -4.4492517e-06, 5.700086e-07, 0.00054767914, -3.7646667e-05, -4.08425e-06, 5.702518e-07, 0.0005280709, -4.0748277e-05, -3.71291e-06, 5.6837143e-07, 0.0005069693, -4.3619326e-05, -3.3367733e-06, 5.644246e-07, 0.00048449088, -4.6254732e-05, -2.957363e-06, 5.584748e-07, 0.00046075453, -4.8650407e-05, -2.576178e-06, 5.505918e-07, 0.00043588094, -5.0803268e-05, -2.194688e-06, 5.4085064e-07, 0.0004099921, -5.271122e-05, -1.8143284e-06, 5.293319e-07, 0.00038321075, -5.4373137e-05, -1.436496e-06, 5.1612096e-07, 0.00035566, -5.5788845e-05, -1.0625445e-06, 5.013074e-07, 0.00032746283, -5.69591e-05, -6.9378035e-07, 4.8498487e-07, 0.00029874156, -5.7885554e-05, -3.3145923e-07, 4.6725037e-07, 0.0002696175, -5.8570742e-05, 2.3217734e-08, 4.4820402e-07, 0.00024021049, -5.9018043e-05, 3.6910714e-07, 4.2794838e-07, 0.00021063843, -5.9231643e-05, 7.051261e-07, 4.065882e-07, 0.00018101699, -5.921651e-05, 1.0302551e-06, 3.8422993e-07, 0.00015145913, -5.897834e-05, 1.3435401e-06, 3.6098115e-07, 0.0001220748, -5.8523547e-05, 1.6440946e-06, 3.3695028e-07, 9.297055e-05, -5.785918e-05, 1.9311012e-06, 3.1224604e-07, 6.4249296e-05, -5.6992914e-05, 2.203814e-06, 2.8697718e-07, 3.6009948e-05, -5.5933e-05, 2.4615574e-06, 2.6125187e-07, 8.347148e-06, -5.4688207e-05, 2.70373e-06, 2.3517745e-07, -1.8648954e-05, -5.326779e-05, 2.9298028e-06, 2.0886e-07, -4.4892953e-05, -5.1681443e-05, 3.13932e-06, 1.8240398e-07, -7.0304384e-05, -4.9939234e-05, 3.331899e-06, 1.5591182e-07, -9.48079e-05, -4.8051577e-05, 3.5072312e-06, 1.2948367e-07, -0.00011833347, -4.602918e-05, 3.665079e-06, 1.03217005e-07, -0.00014081642, -4.3882996e-05, 3.8052772e-06, 7.7206366e-08, -0.00016219766, -4.1624175e-05, 3.9277306e-06, 5.1543033e-08, -0.00018242367, -3.9264014e-05, 4.032413e-06, 2.6314797e-08, -0.00020144664, -3.6813915e-05, 4.119366e-06, 1.6056904e-09, -0.00021922447, -3.4285353e-05, 4.188697e-06, -2.2504235e-08, -0.00023572078, -3.1689793e-05, 4.2405763e-06, -4.593911e-08, -0.00025090497, -2.903869e-05, 4.2752363e-06, -6.8627436e-08, -0.00026475207, -2.6343421e-05, 4.2929682e-06, -9.0502255e-08, -0.00027724289, -2.361525e-05, 4.294121e-06, -1.1150127e-07, -0.00028836366, -2.086529e-05, 4.2790953e-06, -1.3156702e-07, -0.00029810632, -1.8104458e-05, 4.248345e-06, -1.5064691e-07, -0.00030646808, -1.5343456e-05, 4.2023707e-06, -1.6869333e-07, -0.00031345146, -1.2592711e-05, 4.1417193e-06, -1.8566374e-07, -0.00031906416, -9.862363e-06, 4.066978e-06, -2.0152062e-07, -0.00032331882, -7.1622253e-06, 3.9787747e-06, -2.1623163e-07, -0.00032623296, -4.5017537e-06, 3.8777707e-06, -2.2976944e-07, -0.0003278287, -1.890025e-06, 3.7646605e-06, -2.4211184e-07, -0.00032813253, 6.642919e-07, 3.6401673e-06, -2.532417e-07, -0.0003271753, 3.152957e-06, 3.5050389e-06, -2.6314675e-07, -0.00032499182, 5.5681808e-06, 3.3600452e-06, -2.7181972e-07, -0.00032162058, 7.902641e-06, 3.2059747e-06, -2.7925813e-07, -0.00031710375, 1.0149502e-05, 3.0436304e-06, -2.854642e-07, -0.00031148674, 1.2302423e-05, 2.8738268e-06, -2.9044477e-07, -0.00030481795, 1.4355575e-05, 2.6973871e-06, -2.9421102e-07, -0.00029714865, 1.6303653e-05, 2.515139e-06, -2.9677855e-07, -0.0002885326, 1.8141869e-05, 2.3279115e-06, -2.9816704e-07, -0.00027902581, 1.9865978e-05, 2.1365333e-06, -2.984001e-07, -0.00026868627, 2.1472262e-05, 1.9418271e-06, -2.9750515e-07, -0.0002575737, 2.2957545e-05, 1.744609e-06, -2.955132e-07, -0.00024574934, 2.431918e-05, 1.545684e-06, -2.9245857e-07, -0.0002332755, 2.5555057e-05, 1.3458441e-06, -2.8837883e-07, -0.0002202155, 2.6663587e-05, 1.1458654e-06, -2.8331442e-07, -0.00020663331, 2.7643708e-05, 9.4650557e-07, -2.7730857e-07, -0.00019259329, 2.8494866e-05, 7.485012e-07, -2.7040693e-07, -0.00017815996, 2.9217003e-05, 5.5256595e-07, -2.6265744e-07, -0.00016339774, 2.9810557e-05, 3.5938814e-07, -2.5411012e-07, -0.0001483707, 3.0276437e-05, 1.6962883e-07, -2.4481665e-07, -0.00013314236, 3.0616015e-05, -1.6079946e-08, -2.3483035e-07, -0.000117775446, 3.08311e-05, -1.9713693e-07, -2.2420585e-07, -0.00010233165, 3.0923933e-05, -3.7297312e-07, -2.129988e-07, -8.6871456e-05, 3.0897165e-05, -5.430531e-07, -2.0126572e-07, -7.145393e-05, 3.0753825e-05, -7.068763e-07, -1.8906374e-07, -5.6136512e-05, 3.0497315e-05, -8.63978e-07, -1.7645031e-07, -4.097487e-05, 3.0131378e-05, -1.0139303e-06, -1.634831e-07, -2.6022713e-05, 2.9660077e-05, -1.1563425e-06, -1.5021962e-07, -1.1331644e-05, 2.9087783e-05, -1.2908621e-06, -1.3671718e-07, 3.04899e-06, 2.8419128e-05, -1.417175e-06, -1.230325e-07};
	localparam real hb[0:1199] = {0.02089113, 3.3151082e-05, -4.3065935e-05, -1.3363545e-07, 0.020857995, 9.934768e-05, -4.2787167e-05, -3.9975208e-07, 0.020791832, 0.00016522867, -4.223146e-05, -6.624789e-07, 0.020692853, 0.00023058585, -4.1402196e-05, -9.197127e-07, 0.020561367, 0.00029521363, -4.030422e-05, -1.1694873e-06, 0.020397792, 0.00035890998, -3.8943755e-05, -1.4099754e-06, 0.020202644, 0.00042147728, -3.7328326e-05, -1.63949e-06, 0.019976534, 0.0004827232, -3.5466684e-05, -1.8564855e-06, 0.01972017, 0.0005424616, -3.336872e-05, -2.0595573e-06, 0.019434351, 0.0006005129, -3.1045372e-05, -2.247443e-06, 0.019119965, 0.00065670535, -2.850855e-05, -2.4190206e-06, 0.018777981, 0.00071087515, -2.5771038e-05, -2.573307e-06, 0.018409451, 0.0007628674, -2.2846416e-05, -2.7094582e-06, 0.0180155, 0.00081253634, -1.9748964e-05, -2.8267657e-06, 0.017597325, 0.0008597462, -1.649358e-05, -2.9246546e-06, 0.017156184, 0.00090437126, -1.309568e-05, -3.0026804e-06, 0.016693402, 0.0009462965, -9.5711275e-06, -3.0605268e-06, 0.016210355, 0.0009854177, -5.936136e-06, -3.0980007e-06, 0.015708467, 0.0010216419, -2.2071874e-06, -3.1150287e-06, 0.015189208, 0.0010548875, 1.5990514e-06, -3.1116538e-06, 0.014654087, 0.0010850846, 5.465811e-06, -3.0880294e-06, 0.014104641, 0.0011121746, 9.376297e-06, -3.0444157e-06, 0.013542437, 0.001136111, 1.3313769e-05, -2.9811733e-06, 0.012969061, 0.0011568589, 1.7261615e-05, -2.89876e-06, 0.012386113, 0.0011743947, 2.1203417e-05, -2.7977223e-06, 0.011795203, 0.0011887072, 2.5123034e-05, -2.6786931e-06, 0.011197943, 0.0011997957, 2.9004652e-05, -2.5423833e-06, 0.010595943, 0.0012076716, 3.2832853e-05, -2.3895775e-06, 0.009990803, 0.0012123566, 3.659268e-05, -2.221127e-06, 0.009384112, 0.0012138837, 4.0269675e-05, -2.0379443e-06, 0.008777439, 0.0012122962, 4.3849952e-05, -1.8409968e-06, 0.008172326, 0.0012076475, 4.732023e-05, -1.6313006e-06, 0.0075702905, 0.0012000008, 5.0667884e-05, -1.4099147e-06, 0.006972813, 0.0011894285, 5.3880976e-05, -1.1779345e-06, 0.006381336, 0.0011760121, 5.6948305e-05, -9.364856e-07, 0.00579726, 0.0011598415, 5.9859427e-05, -6.867187e-07, 0.0052219373, 0.0011410147, 6.260469e-05, -4.2980258e-07, 0.0046566706, 0.0011196368, 6.5175256e-05, -1.6691912e-07, 0.0041027074, 0.0010958203, 6.7563116e-05, 1.00742795e-07, 0.0035612374, 0.0010696838, 6.976111e-05, 3.7199266e-07, 0.0030333898, 0.0010413518, 7.176296e-05, 6.456437e-07, 0.0025202301, 0.0010109541, 7.356322e-05, 9.2051806e-07, 0.002022758, 0.0009786253, 7.515736e-05, 1.1954519e-06, 0.0015419039, 0.000944504, 7.65417e-05, 1.4693001e-06, 0.0010785293, 0.0009087323, 7.7713434e-05, 1.7409408e-06, 0.00063342287, 0.00087145536, 7.867064e-05, 2.0092798e-06, 0.00020730059, 0.00083282066, 7.941223e-05, 2.273255e-06, -0.000199196, 0.0007929776, 7.993798e-05, 2.531839e-06, -0.0005855002, 0.0007520764, 8.024848e-05, 2.7840447e-06, -0.00095112086, 0.00071026833, 8.034514e-05, 3.028927e-06, -0.0012956422, 0.0006677045, 8.023015e-05, 3.2655869e-06, -0.0016187241, 0.0006245356, 7.990647e-05, 3.493173e-06, -0.0019201015, 0.00058091135, 7.937779e-05, 3.7108857e-06, -0.002199584, 0.0005369799, 7.86485e-05, 3.9179786e-06, -0.002457054, 0.00049288716, 7.772369e-05, 4.1137596e-06, -0.0026924678, 0.00044877693, 7.660907e-05, 4.297595e-06, -0.0029058512, 0.00040478964, 7.5310956e-05, 4.4689077e-06, -0.0030973004, 0.0003610625, 7.383625e-05, 4.6271816e-06, -0.003266979, 0.00031772873, 7.219238e-05, 4.77196e-06, -0.0034151159, 0.00027491737, 7.038726e-05, 4.9028476e-06, -0.0035420037, 0.0002327528, 6.842926e-05, 5.01951e-06, -0.003647996, 0.00019135444, 6.632717e-05, 5.1216743e-06, -0.0037335046, 0.00015083635, 6.409014e-05, 5.209129e-06, -0.003798997, 0.00011130705, 6.172764e-05, 5.281723e-06, -0.0038449934, 7.286914e-05, 5.924944e-05, 5.3393655e-06, -0.003872064, 3.561914e-05, 5.666554e-05, 5.3820245e-06, -0.0038808254, -3.5276486e-07, 5.398614e-05, 5.4097272e-06, -0.003871938, -3.49629e-05, 5.12216e-05, 5.4225566e-06, -0.003846102, -6.813426e-05, 4.8382382e-05, 5.420651e-06, -0.003804055, -9.979662e-05, 4.547903e-05, 5.404204e-06, -0.0037465673, -0.00012988667, 4.2522115e-05, 5.373458e-06, -0.0036744396, -0.00015834805, 3.9522194e-05, 5.3287076e-06, -0.0035884988, -0.00018513142, 3.6489775e-05, 5.270295e-06, -0.003489595, -0.00021019446, 3.343528e-05, 5.198606e-06, -0.003378597, -0.0002335019, 3.0369003e-05, 5.1140705e-06, -0.0032563903, -0.0002550254, 2.7301081e-05, 5.017158e-06, -0.0031238724, -0.00027474365, 2.4241448e-05, 4.908377e-06, -0.00298195, -0.0002926421, 2.1199816e-05, 4.7882686e-06, -0.002831535, -0.00030871294, 1.8185634e-05, 4.657408e-06, -0.002673542, -0.000322955, 1.5208058e-05, 4.5163997e-06, -0.002508884, -0.0003353736, 1.2275935e-05, 4.365872e-06, -0.0023384704, -0.00034598025, 9.39776e-06, 4.2064794e-06, -0.002163203, -0.00035479266, 6.5816644e-06, 4.0388954e-06, -0.001983973, -0.0003618344, 3.83539e-06, 3.863811e-06, -0.0018016589, -0.00036713466, 1.1662675e-06, 3.6819313e-06, -0.0016171229, -0.00037072808, -1.4188005e-06, 3.4939735e-06, -0.0014312087, -0.00037265453, -3.9133556e-06, 3.3006627e-06, -0.0012447389, -0.0003729587, -6.3113976e-06, 3.1027296e-06, -0.0010585124, -0.00037168985, -8.607398e-06, 2.900908e-06, -0.00087330246, -0.00036890176, -1.0796308e-05, 2.6959303e-06, -0.00068985444, -0.00036465205, -1.2873567e-05, 2.4885273e-06, -0.00050888397, -0.00035900212, -1.4835111e-05, 2.2794236e-06, -0.00033107505, -0.00035201685, -1.6677372e-05, 2.0693353e-06, -0.00015707855, -0.00034376408, -1.8397284e-05, 1.8589683e-06, 1.2489361e-05, -0.00033431454, -1.9992282e-05, 1.6490147e-06, 0.0001770485, -0.00032374132, -2.1460299e-05, 1.4401517e-06, 0.0003360557, -0.0003121196, -2.2799763e-05, 1.2330385e-06, 0.000489006, -0.00029952647, -2.4009592e-05, 1.0283145e-06, 0.0006354331, -0.0002860403, -2.508919e-05, 8.265978e-07, 0.00077491056, -0.0002717408, -2.6038428e-05, 6.2848255e-07, 0.00090705155, -0.00025670833, -2.6857646e-05, 4.3453778e-07, 0.00103151, -0.0002410238, -2.7547636e-05, 2.4530576e-07, 0.00114798, -0.00022476834, -2.8109625e-05, 6.130047e-08, 0.0012561965, -0.00020802299, -2.8545266e-05, -1.1699363e-07, 0.0013559345, -0.0001908683, -2.8856623e-05, -2.8912274e-07, 0.0014470097, -0.00017338422, -2.9046143e-05, -4.5466476e-07, 0.0015292768, -0.00015564967, -2.9116654e-05, -6.132301e-07, 0.0016026304, -0.00013774236, -2.9071338e-05, -7.6446247e-07, 0.001667003, -0.00011973852, -2.8913702e-05, -9.080394e-07, 0.0017223652, -0.00010171263, -2.864758e-05, -1.0436728e-06, 0.001768724, -8.37372e-05, -2.8277087e-05, -1.1711089e-06, 0.0018061224, -6.588259e-05, -2.7806615e-05, -1.290129e-06, 0.0018346378, -4.8216738e-05, -2.7240796e-05, -1.400549e-06, 0.0018543813, -3.080503e-05, -2.65845e-05, -1.5022194e-06, 0.0018654956, -1.3710084e-05, -2.5842783e-05, -1.5950253e-06, 0.001868154, 3.008397e-06, -2.502089e-05, -1.6788858e-06, 0.0018625592, 1.9293771e-05, -2.412422e-05, -1.7537535e-06, 0.0018489413, 3.5092595e-05, -2.3158298e-05, -1.8196142e-06, 0.001827556, 5.0354738e-05, -2.2128765e-05, -1.876486e-06, 0.0017986838, 6.503348e-05, -2.1041336e-05, -1.924418e-06, 0.001762627, 7.908561e-05, -1.99018e-05, -1.963491e-06, 0.0017197091, 9.2471484e-05, -1.8715973e-05, -1.9938143e-06, 0.0016702726, 0.000105155086, -1.74897e-05, -2.0155262e-06, 0.0016146766, 0.00011710408, -1.6228809e-05, -2.0287923e-06, 0.0015532956, 0.00012828982, -1.4939109e-05, -2.0338043e-06, 0.0014865181, 0.00013868736, -1.362636e-05, -2.0307787e-06, 0.0014147433, 0.00014827549, -1.2296254e-05, -2.0199554e-06, 0.0013383805, 0.00015703666, -1.0954395e-05, -2.0015964e-06, 0.0012578468, 0.000164957, -9.606287e-06, -1.975984e-06, 0.0011735654, 0.00017202628, -8.257306e-06, -1.9434199e-06, 0.0010859636, 0.00017823778, -6.912691e-06, -1.9042225e-06, 0.0009954711, 0.00018358832, -5.577525e-06, -1.8587268e-06, 0.00090251875, 0.00018807813, -4.2567203e-06, -1.8072818e-06, 0.00080753595, 0.0001917108, -2.955006e-06, -1.750249e-06, 0.00071094977, 0.00019449311, -1.676913e-06, -1.688001e-06, 0.000613183, 0.000196435, -4.2676385e-07, -1.6209199e-06, 0.0005146528, 0.00019754937, 7.913391e-07, -1.5493953e-06, 0.00041576906, 0.00019785204, 1.9735228e-06, -1.4738231e-06, 0.0003169331, 0.00019736159, 3.1161526e-06, -1.3946036e-06, 0.00021853628, 0.00019609914, 4.215839e-06, -1.3121403e-06, 0.000120958815, 0.00019408834, 5.2694445e-06, -1.2268376e-06, 2.4568484e-05, 0.00019135511, 6.27409e-06, -1.1391004e-06, -7.0280425e-05, 0.00018792751, 7.227157e-06, -1.0493314e-06, -0.00016324816, 0.00018383561, 8.1262915e-06, -9.579305e-07, -0.0002540105, 0.00017911129, 8.969408e-06, -8.6529326e-07, -0.00034225947, 0.00017378808, 9.754686e-06, -7.7180914e-07, -0.00042770442, 0.00016790099, 1.0480577e-05, -6.778606e-07, -0.0005100724, 0.00016148636, 1.1145795e-05, -5.838219e-07, -0.00058910897, 0.00015458165, 1.1749322e-05, -4.900576e-07, -0.00066457863, 0.0001472253, 1.22904e-05, -3.9692156e-07, -0.0007362654, 0.00013945656, 1.27685325e-05, -3.047562e-07, -0.00080397294, 0.00013131526, 1.3183473e-05, -2.138912e-07, -0.0008675251, 0.00012284175, 1.3535224e-05, -1.2464257e-07, -0.00092676596, 0.00011407665, 1.3824031e-05, -3.7312006e-08, -0.0009815599, 0.000105060666, 1.4050373e-05, 4.781396e-08, -0.0010317914, 9.583455e-05, 1.4214956e-05, 1.3046464e-07, -0.001077366, 8.643882e-05, 1.4318705e-05, 2.103858e-07, -0.0011182086, 7.691369e-05, 1.4362755e-05, 2.8734019e-07, -0.0011542646, 6.729886e-05, 1.43484385e-05, 3.6110802e-07, -0.0011854989, 5.7633446e-05, 1.427728e-05, 4.3148725e-07, -0.0012118958, 4.7955797e-05, 1.4150984e-05, 4.9829407e-07, -0.0012334588, 3.8303377e-05, 1.3971419e-05, 5.61363e-07, -0.0012502094, 2.8712651e-05, 1.3740616e-05, 6.205469e-07, -0.0012621875, 1.9218973e-05, 1.3460747e-05, 6.7571756e-07, -0.0012694502, 9.856461e-06, 1.31341185e-05, 7.2676505e-07, -0.0012720713, 6.579164e-07, 1.276316e-05, 7.735982e-07, -0.0012701406, -8.345278e-06, 1.2350408e-05, 8.1614405e-07, -0.0012637634, -1.7123242e-05, 1.1898494e-05, 8.543481e-07, -0.0012530595, -2.5647678e-05, 1.1410139e-05, 8.881737e-07, -0.0012381624, -3.389193e-05, 1.0888131e-05, 9.176018e-07, -0.0012192184, -4.1831066e-05, 1.03353195e-05, 9.4263083e-07, -0.0011963861, -4.9441896e-05, 9.7546e-06, 9.632757e-07, -0.0011698348, -5.6703062e-05, 9.148904e-06, 9.795682e-07, -0.0011397444, -6.3595035e-05, 8.521183e-06, 9.915556e-07, -0.0011063041, -7.010016e-05, 7.874404e-06, 9.993003e-07, -0.0010697114, -7.6202705e-05, 7.2115313e-06, 1.0028796e-06, -0.0010301708, -8.1888815e-05, 6.535516e-06, 1.0023847e-06, -0.0009878939, -8.7146575e-05, 5.849289e-06, 9.979202e-07, -0.00094309734, -9.1965965e-05, 5.1557467e-06, 9.89603e-07, -0.0008960024, -9.6338896e-05, 4.457742e-06, 9.775619e-07, -0.0008468339, -0.00010025915, 3.7580744e-06, 9.619366e-07, -0.00079581945, -0.00010372239, 3.0594817e-06, 9.428773e-07, -0.00074318814, -0.000106726126, 2.36463e-06, 9.205432e-07, -0.00068917003, -0.000109269655, 1.6761053e-06, 8.9510223e-07, -0.00063399505, -0.00011135404, 9.964059e-07, 8.6673e-07, -0.00057789206, -0.00011298208, 3.2793542e-07, 8.356088e-07, -0.0005210883, -0.000114158225, -3.2700433e-07, 8.0192706e-07, -0.00046380822, -0.000114888535, -9.662197e-07, 7.658782e-07, -0.00040627285, -0.000115180614, -1.5876305e-06, 7.2765994e-07, -0.00034869916, -0.00011504354, -2.1892758e-06, 6.8747323e-07, -0.00029129916, -0.000114487826, -2.7693175e-06, 6.455217e-07, -0.00023427921, -0.00011352528, -3.3260449e-06, 6.020107e-07, -0.00017783955, -0.000112169015, -3.8578783e-06, 5.571463e-07, -0.00012217351, -0.000110433284, -4.363371e-06, 5.111347e-07, -6.746702e-05, -0.00010833344, -4.841212e-06, 4.6418145e-07, -1.38980895e-05, -0.00010588588, -5.2902283e-06, 4.164905e-07, 3.8363713e-05, -0.00010310789, -5.7093844e-06, 3.682637e-07, 8.915767e-05, -0.00010001759, -6.097784e-06, 3.1969986e-07, 0.00013833233, -9.6633885e-05, -6.4546707e-06, 2.7099426e-07, 0.00018574584, -9.2976305e-05, -6.779425e-06, 2.2233787e-07, 0.00023126627, -8.906495e-05, -7.0715655e-06, 1.7391679e-07, 0.00027477185, -8.492043e-05, -7.330747e-06, 1.2591161e-07, 0.00031615124, -8.0563696e-05, -7.5567577e-06, 7.8496946e-08, 0.00035530367, -7.6016026e-05, -7.749518e-06, 3.1840855e-08, 0.00039213896, -7.129892e-05, -7.909074e-06, -1.38956295e-08, 0.00042657787, -6.643398e-05, -8.035602e-06, -5.855892e-08, 0.00045855186, -6.1442865e-05, -8.129394e-06, -1.020033e-07, 0.00048800325, -5.634719e-05, -8.190864e-06, -1.4409123e-07, 0.0005148851, -5.116844e-05, -8.220535e-06, -1.8469376e-07, 0.0005391613, -4.5927904e-05, -8.219043e-06, -2.236907e-07, 0.0005608062, -4.06466e-05, -8.187122e-06, -2.6097098e-07, 0.00057980453, -3.534518e-05, -8.125607e-06, -2.964327e-07, 0.00059615134, -3.00439e-05, -8.035425e-06, -3.299834e-07, 0.0006098517, -2.4762514e-05, -7.917587e-06, -3.6154026e-07, 0.0006209203, -1.9520232e-05, -7.773189e-06, -3.9102994e-07, 0.00062938145, -1.4335658e-05, -7.603398e-06, -4.183888e-07, 0.0006352685, -9.226734e-06, -7.4094505e-06, -4.4356287e-07, 0.00063862366, -4.210683e-06, -7.192644e-06, -4.6650783e-07, 0.0006394974, 6.9603163e-07, -6.954332e-06, -4.8718886e-07, 0.0006379484, 5.4777533e-06, -6.6959183e-06, -5.055807e-07, 0.0006340429, 1.0119673e-05, -6.4188466e-06, -5.216673e-07, 0.0006278543, 1.460786e-05, -6.1245987e-06, -5.3544187e-07, 0.0006194628, 1.89293e-05, -5.8146848e-06, -5.469065e-07, 0.0006089548, 2.3071916e-05, -5.490638e-06, -5.560721e-07, 0.0005964225, 2.7024593e-05, -5.1540096e-06, -5.62958e-07, 0.00058196357, 3.0777202e-05, -4.806359e-06, -5.6759166e-07, 0.0005656802, 3.43206e-05, -4.4492517e-06, -5.700086e-07, 0.00054767914, 3.7646667e-05, -4.08425e-06, -5.702518e-07, 0.0005280709, 4.0748277e-05, -3.71291e-06, -5.6837143e-07, 0.0005069693, 4.3619326e-05, -3.3367733e-06, -5.644246e-07, 0.00048449088, 4.6254732e-05, -2.957363e-06, -5.584748e-07, 0.00046075453, 4.8650407e-05, -2.576178e-06, -5.505918e-07, 0.00043588094, 5.0803268e-05, -2.194688e-06, -5.4085064e-07, 0.0004099921, 5.271122e-05, -1.8143284e-06, -5.293319e-07, 0.00038321075, 5.4373137e-05, -1.436496e-06, -5.1612096e-07, 0.00035566, 5.5788845e-05, -1.0625445e-06, -5.013074e-07, 0.00032746283, 5.69591e-05, -6.9378035e-07, -4.8498487e-07, 0.00029874156, 5.7885554e-05, -3.3145923e-07, -4.6725037e-07, 0.0002696175, 5.8570742e-05, 2.3217734e-08, -4.4820402e-07, 0.00024021049, 5.9018043e-05, 3.6910714e-07, -4.2794838e-07, 0.00021063843, 5.9231643e-05, 7.051261e-07, -4.065882e-07, 0.00018101699, 5.921651e-05, 1.0302551e-06, -3.8422993e-07, 0.00015145913, 5.897834e-05, 1.3435401e-06, -3.6098115e-07, 0.0001220748, 5.8523547e-05, 1.6440946e-06, -3.3695028e-07, 9.297055e-05, 5.785918e-05, 1.9311012e-06, -3.1224604e-07, 6.4249296e-05, 5.6992914e-05, 2.203814e-06, -2.8697718e-07, 3.6009948e-05, 5.5933e-05, 2.4615574e-06, -2.6125187e-07, 8.347148e-06, 5.4688207e-05, 2.70373e-06, -2.3517745e-07, -1.8648954e-05, 5.326779e-05, 2.9298028e-06, -2.0886e-07, -4.4892953e-05, 5.1681443e-05, 3.13932e-06, -1.8240398e-07, -7.0304384e-05, 4.9939234e-05, 3.331899e-06, -1.5591182e-07, -9.48079e-05, 4.8051577e-05, 3.5072312e-06, -1.2948367e-07, -0.00011833347, 4.602918e-05, 3.665079e-06, -1.03217005e-07, -0.00014081642, 4.3882996e-05, 3.8052772e-06, -7.7206366e-08, -0.00016219766, 4.1624175e-05, 3.9277306e-06, -5.1543033e-08, -0.00018242367, 3.9264014e-05, 4.032413e-06, -2.6314797e-08, -0.00020144664, 3.6813915e-05, 4.119366e-06, -1.6056904e-09, -0.00021922447, 3.4285353e-05, 4.188697e-06, 2.2504235e-08, -0.00023572078, 3.1689793e-05, 4.2405763e-06, 4.593911e-08, -0.00025090497, 2.903869e-05, 4.2752363e-06, 6.8627436e-08, -0.00026475207, 2.6343421e-05, 4.2929682e-06, 9.0502255e-08, -0.00027724289, 2.361525e-05, 4.294121e-06, 1.1150127e-07, -0.00028836366, 2.086529e-05, 4.2790953e-06, 1.3156702e-07, -0.00029810632, 1.8104458e-05, 4.248345e-06, 1.5064691e-07, -0.00030646808, 1.5343456e-05, 4.2023707e-06, 1.6869333e-07, -0.00031345146, 1.2592711e-05, 4.1417193e-06, 1.8566374e-07, -0.00031906416, 9.862363e-06, 4.066978e-06, 2.0152062e-07, -0.00032331882, 7.1622253e-06, 3.9787747e-06, 2.1623163e-07, -0.00032623296, 4.5017537e-06, 3.8777707e-06, 2.2976944e-07, -0.0003278287, 1.890025e-06, 3.7646605e-06, 2.4211184e-07, -0.00032813253, -6.642919e-07, 3.6401673e-06, 2.532417e-07, -0.0003271753, -3.152957e-06, 3.5050389e-06, 2.6314675e-07, -0.00032499182, -5.5681808e-06, 3.3600452e-06, 2.7181972e-07, -0.00032162058, -7.902641e-06, 3.2059747e-06, 2.7925813e-07, -0.00031710375, -1.0149502e-05, 3.0436304e-06, 2.854642e-07, -0.00031148674, -1.2302423e-05, 2.8738268e-06, 2.9044477e-07, -0.00030481795, -1.4355575e-05, 2.6973871e-06, 2.9421102e-07, -0.00029714865, -1.6303653e-05, 2.515139e-06, 2.9677855e-07, -0.0002885326, -1.8141869e-05, 2.3279115e-06, 2.9816704e-07, -0.00027902581, -1.9865978e-05, 2.1365333e-06, 2.984001e-07, -0.00026868627, -2.1472262e-05, 1.9418271e-06, 2.9750515e-07, -0.0002575737, -2.2957545e-05, 1.744609e-06, 2.955132e-07, -0.00024574934, -2.431918e-05, 1.545684e-06, 2.9245857e-07, -0.0002332755, -2.5555057e-05, 1.3458441e-06, 2.8837883e-07, -0.0002202155, -2.6663587e-05, 1.1458654e-06, 2.8331442e-07, -0.00020663331, -2.7643708e-05, 9.4650557e-07, 2.7730857e-07, -0.00019259329, -2.8494866e-05, 7.485012e-07, 2.7040693e-07, -0.00017815996, -2.9217003e-05, 5.5256595e-07, 2.6265744e-07, -0.00016339774, -2.9810557e-05, 3.5938814e-07, 2.5411012e-07, -0.0001483707, -3.0276437e-05, 1.6962883e-07, 2.4481665e-07, -0.00013314236, -3.0616015e-05, -1.6079946e-08, 2.3483035e-07, -0.000117775446, -3.08311e-05, -1.9713693e-07, 2.2420585e-07, -0.00010233165, -3.0923933e-05, -3.7297312e-07, 2.129988e-07, -8.6871456e-05, -3.0897165e-05, -5.430531e-07, 2.0126572e-07, -7.145393e-05, -3.0753825e-05, -7.068763e-07, 1.8906374e-07, -5.6136512e-05, -3.0497315e-05, -8.63978e-07, 1.7645031e-07, -4.097487e-05, -3.0131378e-05, -1.0139303e-06, 1.634831e-07, -2.6022713e-05, -2.9660077e-05, -1.1563425e-06, 1.5021962e-07, -1.1331644e-05, -2.9087783e-05, -1.2908621e-06, 1.3671718e-07, 3.04899e-06, -2.8419128e-05, -1.417175e-06, 1.230325e-07};
endpackage
`endif
