`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam N = 4;
	localparam real Lfr[0:3] = {0.98584217, 0.98584217, 0.9781171, 0.9781171};
	localparam real Lfi[0:3] = {0.10665247, -0.10665247, 0.041062612, -0.041062612};
	localparam real Lbr[0:3] = {0.98584217, 0.98584217, 0.9781171, 0.9781171};
	localparam real Lbi[0:3] = {0.10665247, -0.10665247, 0.041062612, -0.041062612};
	localparam real Wfr[0:3] = {8.595155e-05, 8.595155e-05, -2.8021776e-05, -2.8021776e-05};
	localparam real Wfi[0:3] = {0.00010408412, -0.00010408412, -0.00011768973, 0.00011768973};
	localparam real Wbr[0:3] = {-8.595155e-05, -8.595155e-05, 2.8021776e-05, 2.8021776e-05};
	localparam real Wbi[0:3] = {-0.00010408412, 0.00010408412, 0.00011768973, -0.00011768973};
	localparam real Ffr[0:3][0:79] = '{
		'{9.517404, 5.803959, -0.47750285, -0.05147556, 12.334175, 5.4531856, -0.54906327, -0.04322708, 14.961022, 5.045163, -0.61307025, -0.034616325, 17.370718, 4.5855722, -0.66890925, -0.025749026, 19.539005, 4.0805964, -0.7160708, -0.01673212, 21.444826, 3.5368402, -0.75415415, -0.0076724873, 23.070515, 2.9612474, -0.7828705, 0.0013242945, 24.401941, 2.3610132, -0.80204415, 0.010155137, 25.428623, 1.7434981, -0.8116131, 0.018720599, 26.143776, 1.1161392, -0.81162727, 0.026925975, 26.544338, 0.48636296, -0.80224645, 0.034682315, 26.630938, -0.13850014, -0.78373647, 0.041907355, 26.407831, -0.75129956, -0.75646454, 0.04852636, 25.882782, -1.3451439, -0.72089285, 0.054472856, 25.066925, -1.9134767, -0.67757225, 0.059689272, 23.974571, -2.4501464, -0.6271338, 0.064127445, 22.622993, -2.9494712, -0.5702805, 0.06774904, 21.032177, -3.4062963, -0.5077778, 0.07052579, 19.224539, -3.8160453, -0.4404439, 0.07243971, 17.224634, -4.174763, -0.36913893, 0.07348309},
		'{9.517404, 5.803959, -0.47750285, -0.05147556, 12.334175, 5.4531856, -0.54906327, -0.04322708, 14.961022, 5.045163, -0.61307025, -0.034616325, 17.370718, 4.5855722, -0.66890925, -0.025749026, 19.539005, 4.0805964, -0.7160708, -0.01673212, 21.444826, 3.5368402, -0.75415415, -0.0076724873, 23.070515, 2.9612474, -0.7828705, 0.0013242945, 24.401941, 2.3610132, -0.80204415, 0.010155137, 25.428623, 1.7434981, -0.8116131, 0.018720599, 26.143776, 1.1161392, -0.81162727, 0.026925975, 26.544338, 0.48636296, -0.80224645, 0.034682315, 26.630938, -0.13850014, -0.78373647, 0.041907355, 26.407831, -0.75129956, -0.75646454, 0.04852636, 25.882782, -1.3451439, -0.72089285, 0.054472856, 25.066925, -1.9134767, -0.67757225, 0.059689272, 23.974571, -2.4501464, -0.6271338, 0.064127445, 22.622993, -2.9494712, -0.5702805, 0.06774904, 21.032177, -3.4062963, -0.5077778, 0.07052579, 19.224539, -3.8160453, -0.4404439, 0.07243971, 17.224634, -4.174763, -0.36913893, 0.07348309},
		'{-9.3133135, -5.688954, 0.4059951, -0.19382812, -12.087016, -5.4058576, 0.3589503, -0.1867144, -14.719161, -5.122835, 0.31308547, -0.17949237, -17.20994, -4.8404956, 0.2684508, -0.17218217, -19.559843, -4.5594215, 0.2250918, -0.16480333, -21.769638, -4.2801695, 0.18304923, -0.15737464, -23.840376, -4.0032682, 0.14235936, -0.14991428, -25.773354, -3.729219, 0.10305402, -0.14243971, -27.570118, -3.4584966, 0.06516069, -0.1349677, -29.232447, -3.1915488, 0.028702687, -0.12751433, -30.762333, -2.9287965, -0.0063007767, -0.12009496, -32.161976, -2.6706343, -0.03983443, -0.11272424, -33.433758, -2.4174297, -0.071886815, -0.1054161, -34.580254, -2.169525, -0.10245016, -0.09818375, -35.604183, -1.9272362, -0.13152024, -0.09103971, -36.50844, -1.6908544, -0.15909624, -0.08399577, -37.296032, -1.4606457, -0.18518062, -0.077063, -37.970116, -1.2368513, -0.20977895, -0.07025181, -38.533955, -1.0196893, -0.2328998, -0.06357187, -38.990906, -0.8093538, -0.25455457, -0.057032187},
		'{-9.3133135, -5.688954, 0.4059951, -0.19382812, -12.087016, -5.4058576, 0.3589503, -0.1867144, -14.719161, -5.122835, 0.31308547, -0.17949237, -17.20994, -4.8404956, 0.2684508, -0.17218217, -19.559843, -4.5594215, 0.2250918, -0.16480333, -21.769638, -4.2801695, 0.18304923, -0.15737464, -23.840376, -4.0032682, 0.14235936, -0.14991428, -25.773354, -3.729219, 0.10305402, -0.14243971, -27.570118, -3.4584966, 0.06516069, -0.1349677, -29.232447, -3.1915488, 0.028702687, -0.12751433, -30.762333, -2.9287965, -0.0063007767, -0.12009496, -32.161976, -2.6706343, -0.03983443, -0.11272424, -33.433758, -2.4174297, -0.071886815, -0.1054161, -34.580254, -2.169525, -0.10245016, -0.09818375, -35.604183, -1.9272362, -0.13152024, -0.09103971, -36.50844, -1.6908544, -0.15909624, -0.08399577, -37.296032, -1.4606457, -0.18518062, -0.077063, -37.970116, -1.2368513, -0.20977895, -0.07025181, -38.533955, -1.0196893, -0.2328998, -0.06357187, -38.990906, -0.8093538, -0.25455457, -0.057032187}};
	localparam real Ffi[0:3][0:79] = '{
		'{-27.674166, 2.5184734, 0.7343557, -0.07050651, -26.267303, 3.1018236, 0.6730319, -0.07499829, -24.579945, 3.6395042, 0.6049443, -0.07854675, -22.636314, 4.1260557, 0.5309941, -0.08112661, -20.463203, 4.556702, 0.45213553, -0.08272423, -18.089605, 4.927395, 0.36936355, -0.08333755, -15.546351, 5.234846, 0.28370175, -0.08297596, -12.865721, 5.4765563, 0.19619007, -0.08165996, -10.081042, 5.650828, 0.10787244, -0.07942076, -7.2262907, 5.7567725, 0.01978466, -0.076299734, -4.335684, 5.794308, -0.0670575, -0.07234777, -1.4432806, 5.764145, -0.15166967, -0.067624524, 1.4174085, 5.6677656, -0.23310979, -0.062197585, 4.2138014, 5.507394, -0.31048825, -0.056141544, 6.9146056, 5.2859583, -0.38297743, -0.049537037, 9.490159, 5.0070434, -0.44982, -0.042469688, 11.912745, 4.67484, -0.5103369, -0.035029057, 14.156885, 4.294086, -0.56393343, -0.02730752, 16.199587, 3.870001, -0.6101051, -0.019399153, 18.02058, 3.4082193, -0.64844173, -0.011398629},
		'{27.674166, -2.5184734, -0.7343557, 0.07050651, 26.267303, -3.1018236, -0.6730319, 0.07499829, 24.579945, -3.6395042, -0.6049443, 0.07854675, 22.636314, -4.1260557, -0.5309941, 0.08112661, 20.463203, -4.556702, -0.45213553, 0.08272423, 18.089605, -4.927395, -0.36936355, 0.08333755, 15.546351, -5.234846, -0.28370175, 0.08297596, 12.865721, -5.4765563, -0.19619007, 0.08165996, 10.081042, -5.650828, -0.10787244, 0.07942076, 7.2262907, -5.7567725, -0.01978466, 0.076299734, 4.335684, -5.794308, 0.0670575, 0.07234777, 1.4432806, -5.764145, 0.15166967, 0.067624524, -1.4174085, -5.6677656, 0.23310979, 0.062197585, -4.2138014, -5.507394, 0.31048825, 0.056141544, -6.9146056, -5.2859583, 0.38297743, 0.049537037, -9.490159, -5.0070434, 0.44982, 0.042469688, -11.912745, -4.67484, 0.5103369, 0.035029057, -14.156885, -4.294086, 0.56393343, 0.02730752, -16.199587, -3.870001, 0.6101051, 0.019399153, -18.02058, -3.4082193, 0.64844173, 0.011398629},
		'{72.51132, -3.862523, 0.92932385, -0.069947086, 70.54214, -4.0116034, 0.92565876, -0.07637553, 68.502144, -4.1457963, 0.9201421, -0.08237119, 66.39871, -4.2654314, 0.91286284, -0.0879391, 64.23903, -4.370855, 0.90391004, -0.09308498, 62.030117, -4.46243, 0.8933728, -0.097815275, 59.7788, -4.540534, 0.88133967, -0.10213701, 57.491722, -4.6055584, 0.86789906, -0.10605783, 55.175316, -4.657907, 0.85313857, -0.10958592, 52.83582, -4.6979938, 0.83714515, -0.11272999, 50.479256, -4.726241, 0.8200046, -0.115499206, 48.111443, -4.7430816, 0.8018018, -0.117903166, 45.737972, -4.7489524, 0.7826203, -0.11995185, 43.364216, -4.7442975, 0.7625425, -0.12165562, 40.995327, -4.729565, 0.741649, -0.12302513, 38.636227, -4.705206, 0.720019, -0.12407131, 36.291626, -4.6716733, 0.69773, -0.12480536, 33.965984, -4.6294217, 0.6748577, -0.12523866, 31.66356, -4.5789046, 0.6514757, -0.12538281, 29.388365, -4.520576, 0.6276561, -0.12524949},
		'{-72.51132, 3.862523, -0.92932385, 0.069947086, -70.54214, 4.0116034, -0.92565876, 0.07637553, -68.502144, 4.1457963, -0.9201421, 0.08237119, -66.39871, 4.2654314, -0.91286284, 0.0879391, -64.23903, 4.370855, -0.90391004, 0.09308498, -62.030117, 4.46243, -0.8933728, 0.097815275, -59.7788, 4.540534, -0.88133967, 0.10213701, -57.491722, 4.6055584, -0.86789906, 0.10605783, -55.175316, 4.657907, -0.85313857, 0.10958592, -52.83582, 4.6979938, -0.83714515, 0.11272999, -50.479256, 4.726241, -0.8200046, 0.115499206, -48.111443, 4.7430816, -0.8018018, 0.117903166, -45.737972, 4.7489524, -0.7826203, 0.11995185, -43.364216, 4.7442975, -0.7625425, 0.12165562, -40.995327, 4.729565, -0.741649, 0.12302513, -38.636227, 4.705206, -0.720019, 0.12407131, -36.291626, 4.6716733, -0.69773, 0.12480536, -33.965984, 4.6294217, -0.6748577, 0.12523866, -31.66356, 4.5789046, -0.6514757, 0.12538281, -29.388365, 4.520576, -0.6276561, 0.12524949}};
	localparam real Fbr[0:3][0:79] = '{
		'{-9.517404, 5.803959, 0.47750285, -0.05147556, -12.334175, 5.4531856, 0.54906327, -0.04322708, -14.961022, 5.045163, 0.61307025, -0.034616325, -17.370718, 4.5855722, 0.66890925, -0.025749026, -19.539005, 4.0805964, 0.7160708, -0.01673212, -21.444826, 3.5368402, 0.75415415, -0.0076724873, -23.070515, 2.9612474, 0.7828705, 0.0013242945, -24.401941, 2.3610132, 0.80204415, 0.010155137, -25.428623, 1.7434981, 0.8116131, 0.018720599, -26.143776, 1.1161392, 0.81162727, 0.026925975, -26.544338, 0.48636296, 0.80224645, 0.034682315, -26.630938, -0.13850014, 0.78373647, 0.041907355, -26.407831, -0.75129956, 0.75646454, 0.04852636, -25.882782, -1.3451439, 0.72089285, 0.054472856, -25.066925, -1.9134767, 0.67757225, 0.059689272, -23.974571, -2.4501464, 0.6271338, 0.064127445, -22.622993, -2.9494712, 0.5702805, 0.06774904, -21.032177, -3.4062963, 0.5077778, 0.07052579, -19.224539, -3.8160453, 0.4404439, 0.07243971, -17.224634, -4.174763, 0.36913893, 0.07348309},
		'{-9.517404, 5.803959, 0.47750285, -0.05147556, -12.334175, 5.4531856, 0.54906327, -0.04322708, -14.961022, 5.045163, 0.61307025, -0.034616325, -17.370718, 4.5855722, 0.66890925, -0.025749026, -19.539005, 4.0805964, 0.7160708, -0.01673212, -21.444826, 3.5368402, 0.75415415, -0.0076724873, -23.070515, 2.9612474, 0.7828705, 0.0013242945, -24.401941, 2.3610132, 0.80204415, 0.010155137, -25.428623, 1.7434981, 0.8116131, 0.018720599, -26.143776, 1.1161392, 0.81162727, 0.026925975, -26.544338, 0.48636296, 0.80224645, 0.034682315, -26.630938, -0.13850014, 0.78373647, 0.041907355, -26.407831, -0.75129956, 0.75646454, 0.04852636, -25.882782, -1.3451439, 0.72089285, 0.054472856, -25.066925, -1.9134767, 0.67757225, 0.059689272, -23.974571, -2.4501464, 0.6271338, 0.064127445, -22.622993, -2.9494712, 0.5702805, 0.06774904, -21.032177, -3.4062963, 0.5077778, 0.07052579, -19.224539, -3.8160453, 0.4404439, 0.07243971, -17.224634, -4.174763, 0.36913893, 0.07348309},
		'{9.3133135, -5.688954, -0.4059951, -0.19382812, 12.087016, -5.4058576, -0.3589503, -0.1867144, 14.719161, -5.122835, -0.31308547, -0.17949237, 17.20994, -4.8404956, -0.2684508, -0.17218217, 19.559843, -4.5594215, -0.2250918, -0.16480333, 21.769638, -4.2801695, -0.18304923, -0.15737464, 23.840376, -4.0032682, -0.14235936, -0.14991428, 25.773354, -3.729219, -0.10305402, -0.14243971, 27.570118, -3.4584966, -0.06516069, -0.1349677, 29.232447, -3.1915488, -0.028702687, -0.12751433, 30.762333, -2.9287965, 0.0063007767, -0.12009496, 32.161976, -2.6706343, 0.03983443, -0.11272424, 33.433758, -2.4174297, 0.071886815, -0.1054161, 34.580254, -2.169525, 0.10245016, -0.09818375, 35.604183, -1.9272362, 0.13152024, -0.09103971, 36.50844, -1.6908544, 0.15909624, -0.08399577, 37.296032, -1.4606457, 0.18518062, -0.077063, 37.970116, -1.2368513, 0.20977895, -0.07025181, 38.533955, -1.0196893, 0.2328998, -0.06357187, 38.990906, -0.8093538, 0.25455457, -0.057032187},
		'{9.3133135, -5.688954, -0.4059951, -0.19382812, 12.087016, -5.4058576, -0.3589503, -0.1867144, 14.719161, -5.122835, -0.31308547, -0.17949237, 17.20994, -4.8404956, -0.2684508, -0.17218217, 19.559843, -4.5594215, -0.2250918, -0.16480333, 21.769638, -4.2801695, -0.18304923, -0.15737464, 23.840376, -4.0032682, -0.14235936, -0.14991428, 25.773354, -3.729219, -0.10305402, -0.14243971, 27.570118, -3.4584966, -0.06516069, -0.1349677, 29.232447, -3.1915488, -0.028702687, -0.12751433, 30.762333, -2.9287965, 0.0063007767, -0.12009496, 32.161976, -2.6706343, 0.03983443, -0.11272424, 33.433758, -2.4174297, 0.071886815, -0.1054161, 34.580254, -2.169525, 0.10245016, -0.09818375, 35.604183, -1.9272362, 0.13152024, -0.09103971, 36.50844, -1.6908544, 0.15909624, -0.08399577, 37.296032, -1.4606457, 0.18518062, -0.077063, 37.970116, -1.2368513, 0.20977895, -0.07025181, 38.533955, -1.0196893, 0.2328998, -0.06357187, 38.990906, -0.8093538, 0.25455457, -0.057032187}};
	localparam real Fbi[0:3][0:79] = '{
		'{27.674166, 2.5184734, -0.7343557, -0.07050651, 26.267303, 3.1018236, -0.6730319, -0.07499829, 24.579945, 3.6395042, -0.6049443, -0.07854675, 22.636314, 4.1260557, -0.5309941, -0.08112661, 20.463203, 4.556702, -0.45213553, -0.08272423, 18.089605, 4.927395, -0.36936355, -0.08333755, 15.546351, 5.234846, -0.28370175, -0.08297596, 12.865721, 5.4765563, -0.19619007, -0.08165996, 10.081042, 5.650828, -0.10787244, -0.07942076, 7.2262907, 5.7567725, -0.01978466, -0.076299734, 4.335684, 5.794308, 0.0670575, -0.07234777, 1.4432806, 5.764145, 0.15166967, -0.067624524, -1.4174085, 5.6677656, 0.23310979, -0.062197585, -4.2138014, 5.507394, 0.31048825, -0.056141544, -6.9146056, 5.2859583, 0.38297743, -0.049537037, -9.490159, 5.0070434, 0.44982, -0.042469688, -11.912745, 4.67484, 0.5103369, -0.035029057, -14.156885, 4.294086, 0.56393343, -0.02730752, -16.199587, 3.870001, 0.6101051, -0.019399153, -18.02058, 3.4082193, 0.64844173, -0.011398629},
		'{-27.674166, -2.5184734, 0.7343557, 0.07050651, -26.267303, -3.1018236, 0.6730319, 0.07499829, -24.579945, -3.6395042, 0.6049443, 0.07854675, -22.636314, -4.1260557, 0.5309941, 0.08112661, -20.463203, -4.556702, 0.45213553, 0.08272423, -18.089605, -4.927395, 0.36936355, 0.08333755, -15.546351, -5.234846, 0.28370175, 0.08297596, -12.865721, -5.4765563, 0.19619007, 0.08165996, -10.081042, -5.650828, 0.10787244, 0.07942076, -7.2262907, -5.7567725, 0.01978466, 0.076299734, -4.335684, -5.794308, -0.0670575, 0.07234777, -1.4432806, -5.764145, -0.15166967, 0.067624524, 1.4174085, -5.6677656, -0.23310979, 0.062197585, 4.2138014, -5.507394, -0.31048825, 0.056141544, 6.9146056, -5.2859583, -0.38297743, 0.049537037, 9.490159, -5.0070434, -0.44982, 0.042469688, 11.912745, -4.67484, -0.5103369, 0.035029057, 14.156885, -4.294086, -0.56393343, 0.02730752, 16.199587, -3.870001, -0.6101051, 0.019399153, 18.02058, -3.4082193, -0.64844173, 0.011398629},
		'{-72.51132, -3.862523, -0.92932385, -0.069947086, -70.54214, -4.0116034, -0.92565876, -0.07637553, -68.502144, -4.1457963, -0.9201421, -0.08237119, -66.39871, -4.2654314, -0.91286284, -0.0879391, -64.23903, -4.370855, -0.90391004, -0.09308498, -62.030117, -4.46243, -0.8933728, -0.097815275, -59.7788, -4.540534, -0.88133967, -0.10213701, -57.491722, -4.6055584, -0.86789906, -0.10605783, -55.175316, -4.657907, -0.85313857, -0.10958592, -52.83582, -4.6979938, -0.83714515, -0.11272999, -50.479256, -4.726241, -0.8200046, -0.115499206, -48.111443, -4.7430816, -0.8018018, -0.117903166, -45.737972, -4.7489524, -0.7826203, -0.11995185, -43.364216, -4.7442975, -0.7625425, -0.12165562, -40.995327, -4.729565, -0.741649, -0.12302513, -38.636227, -4.705206, -0.720019, -0.12407131, -36.291626, -4.6716733, -0.69773, -0.12480536, -33.965984, -4.6294217, -0.6748577, -0.12523866, -31.66356, -4.5789046, -0.6514757, -0.12538281, -29.388365, -4.520576, -0.6276561, -0.12524949},
		'{72.51132, 3.862523, 0.92932385, 0.069947086, 70.54214, 4.0116034, 0.92565876, 0.07637553, 68.502144, 4.1457963, 0.9201421, 0.08237119, 66.39871, 4.2654314, 0.91286284, 0.0879391, 64.23903, 4.370855, 0.90391004, 0.09308498, 62.030117, 4.46243, 0.8933728, 0.097815275, 59.7788, 4.540534, 0.88133967, 0.10213701, 57.491722, 4.6055584, 0.86789906, 0.10605783, 55.175316, 4.657907, 0.85313857, 0.10958592, 52.83582, 4.6979938, 0.83714515, 0.11272999, 50.479256, 4.726241, 0.8200046, 0.115499206, 48.111443, 4.7430816, 0.8018018, 0.117903166, 45.737972, 4.7489524, 0.7826203, 0.11995185, 43.364216, 4.7442975, 0.7625425, 0.12165562, 40.995327, 4.729565, 0.741649, 0.12302513, 38.636227, 4.705206, 0.720019, 0.12407131, 36.291626, 4.6716733, 0.69773, 0.12480536, 33.965984, 4.6294217, 0.6748577, 0.12523866, 31.66356, 4.5789046, 0.6514757, 0.12538281, 29.388365, 4.520576, 0.6276561, 0.12524949}};
	localparam real hf[0:1999] = {0.024986578, -0.000116877105, -3.896343e-05, 2.2712003e-07, 0.024869869, -0.0003495672, -3.6725352e-05, 6.683011e-07, 0.02463752, -0.00057908345, -3.2282736e-05, 1.071189e-06, 0.02429164, -0.00080335606, -2.5699466e-05, 1.4122909e-06, 0.023835355, -0.0010203768, -1.7068134e-05, 1.6701244e-06, 0.023272775, -0.0012282217, -6.508329e-06, 1.825436e-06, 0.02260895, -0.0014250721, 5.835373e-06, 1.8613864e-06, 0.021849804, -0.0016092348, 1.979567e-05, 1.7637041e-06, 0.021002075, -0.0017791594, 3.5185032e-05, 1.5208042e-06, 0.020073237, -0.0019334549, 5.1798383e-05, 1.1238726e-06, 0.019071415, -0.0020709035, 6.941594e-05, 5.669145e-07, 0.018005302, -0.0021904726, 8.7806206e-05, -1.5323168e-07, 0.016884053, -0.0022913238, 0.000106729, -1.0369153e-06, 0.015717195, -0.0023728213, 0.00012593858, -2.0817276e-06, 0.014514523, -0.0024345345, 0.00014518676, -3.2825897e-06, 0.01328599, -0.0024762424, 0.000164226, -4.6318687e-06, 0.012041612, -0.0024979326, 0.00018281244, -6.119525e-06, 0.010791358, -0.0024997983, 0.00020070883, -7.733287e-06, 0.009545049, -0.0024822343, 0.00021768737, -9.458844e-06, 0.008312262, -0.0024458296, 0.00023353235, -1.1280068e-05, 0.0071022296, -0.0023913574, 0.00024804258, -1.31792485e-05, 0.0059237573, -0.0023197657, 0.0002610337, -1.5137347e-05, 0.004785133, -0.0022321627, 0.00027234023, -1.7134254e-05, 0.003694055, -0.002129803, 0.00028181716, -1.9149073e-05, 0.0026575602, -0.0020140712, 0.0002893417, -2.116038e-05, 0.0016819648, -0.0018864649, 0.00029481426, -2.3146522e-05, 0.0007728115, -0.0017485761, 0.00029815955, -2.5085883e-05, -6.517271e-05, -0.0016020724, 0.00029932705, -2.6957157e-05, -0.0008281093, -0.0014486772, 0.0002982914, -2.8739623e-05, -0.0015129913, -0.0012901495, 0.00029505236, -3.0413386e-05, -0.002117696, -0.0011282647, 0.0002896347, -3.195963e-05, -0.0026409882, -0.00096479343, 0.0002820874, -3.3360822e-05, -0.003082513, -0.00080148317, 0.00027248287, -3.4600955e-05, -0.0034427792, -0.00064003846, 0.000260916, -3.5665686e-05, -0.0037231334, -0.0004821034, 0.00024750258, -3.6542533e-05, -0.003925726, -0.00032924407, 0.00023237792, -3.7221005e-05, -0.004053466, -0.00018293266, 0.00021569492, -3.76927e-05, -0.0041099745, -4.453296e-05, 0.00019762217, -3.79514e-05, -0.0040995227, 8.471297e-05, 0.00017834186, -3.7993144e-05, -0.0040269704, 0.00020369625, 0.00015804752, -3.7816237e-05, -0.0038976963, 0.00031145103, 0.00013694167, -3.742127e-05, -0.0037175252, 0.00040716256, 0.00011523339, -3.6811085e-05, -0.0034926496, 0.0004901733, 9.3135954e-05, -3.599074e-05, -0.0032295508, 0.00055998715, 7.086427e-05, -3.4967423e-05, -0.002934917, 0.0006162719, 4.8632493e-05, -3.3750366e-05, -0.0026155617, 0.0006588598, 2.6651622e-05, -3.235072e-05, -0.0022783414, 0.0006877456, 5.1271536e-06, -3.0781408e-05, -0.0019300748, 0.00070308376, -1.5743133e-05, -2.9056979e-05, -0.0015774649, 0.0007051833, -3.577129e-05, -2.7193415e-05, -0.0012270228, 0.00069450086, -5.4781158e-05, -2.5207955e-05, -0.00088499615, 0.00067163265, -7.261017e-05, -2.311889e-05, -0.00055730145, 0.0006373044, -8.911096e-05, -2.0945343e-05, -0.0002494623, 0.00059236056, -0.00010415277, -1.8707058e-05, 3.3447053e-05, 0.00053775206, -0.00011762269, -1.6424181e-05, 0.00028685166, 0.00047452268, -0.00012942658, -1.4117025e-05, 0.0005067189, 0.00040379557, -0.0001394899, -1.1805854e-05, 0.00068959437, 0.00032675808, -0.00014775814, -9.510665e-06, 0.0008326304, 0.00024464677, -0.00015419716, -7.2509692e-06, 0.0009336064, 0.00015873181, -0.00015879319, -5.0455933e-06, 0.0009909424, 7.03015e-05, -0.0001615527, -2.9124817e-06, 0.0010037036, -1.9353303e-05, -0.00016250192, -8.6851696e-07, 0.000971598, -0.00010895448, -0.00016168621, 1.0706473e-06, 0.00089496677, -0.00019725144, -0.00015916926, 2.890736e-06, 0.0007747661, -0.0002830354, -0.00015503199, 4.578985e-06, 0.0006125435, -0.0003651528, -0.0001493714, 6.1242554e-06, 0.00041040673, -0.00044251818, -0.00014229909, 7.517124e-06, 0.00017098685, -0.0005141254, -0.00013393987, 8.749958e-06, -0.000102604055, -0.0005790583, -0.00012442996, 9.816967e-06, -0.00040682033, -0.00063650013, -0.00011391535, 1.0714228e-05, -0.0007377343, -0.00068574096, -0.000102549915, 1.1439698e-05, -0.0010910918, -0.00072618475, -9.049353e-05, 1.1993197e-05, -0.0014623696, -0.0007573539, -7.791015e-05, 1.237638e-05, -0.0018468365, -0.0007788933, -6.496585e-05, 1.2592673e-05, -0.002239615, -0.0007905721, -5.1826923e-05, 1.2647208e-05, -0.0026357428, -0.0007922844, -3.8657945e-05, 1.2546729e-05, -0.0030302363, -0.00078404846, -2.5619947e-05, 1.22994825e-05, -0.0034181513, -0.0007660045, -1.2868641e-05, 1.1915097e-05, -0.0037946438, -0.0007384107, -5.527264e-07, 1.1404446e-05, -0.0041550267, -0.00070163846, 1.1187671e-05, 1.0779499e-05, -0.0044948263, -0.000656166, 2.2222448e-05, 1.0053163e-05, -0.004809833, -0.00060257106, 3.2432832e-05, 9.239121e-06, -0.005096149, -0.0005415224, 4.1712527e-05, 8.351654e-06, -0.0053502326, -0.00047377063, 4.9968694e-05, 7.4054738e-06, -0.0055689337, -0.0004001377, 5.7122783e-05, 6.415538e-06, -0.005749531, -0.00032150644, 6.311115e-05, 5.3968797e-06, -0.005889757, -0.00023880896, 6.788551e-05, 4.3644327e-06, -0.005987819, -0.00015301503, 7.1413204e-05, 3.33286e-06, -0.0060424167, -6.5120075e-05, 7.367729e-05, 2.3163923e-06, -0.0060527516, 2.3866987e-05, 7.467643e-05, 1.3286729e-06, -0.006018531, 0.00011293571, 7.442458e-05, 3.8261123e-07, -0.0059399647, 0.00020108608, 7.295059e-05, -5.097503e-07, -0.005817757, 0.00028734, 7.029756e-05, -1.3373586e-06, -0.0056530945, 0.00037075247, 6.652203e-05, -2.0902578e-06, -0.005447625, 0.00045042214, 6.169313e-05, -2.759682e-06, -0.0052034347, 0.00052550115, 5.589148e-05, -3.3381343e-06, -0.004923017, 0.00059520424, 4.9208058e-05, -3.819447e-06, -0.004609243, 0.00065881707, 4.1742933e-05, -4.198827e-06, -0.0042653196, 0.0007157032, 3.3603916e-05, -4.472884e-06, -0.003894752, 0.0007653107, 2.4905143e-05, -4.639643e-06, -0.0035012984, 0.0008071772, 1.5765636e-05, -4.698537e-06, -0.003088926, 0.0008409337, 6.307793e-06, -4.6503856e-06, -0.0026617618, 0.0008663077, -3.3441117e-06, -4.4973604e-06, -0.0022240446, 0.00088312494, -1.3065424e-05, -4.2429283e-06, -0.0017800763, 0.0008913099, -2.2732595e-05, -3.8917874e-06, -0.0013341709, 0.000890885, -3.2224616e-05, -3.4497868e-06, -0.0008906079, 0.00088196935, -4.142441e-05, -2.9238345e-06, -0.0004535831, 0.00086477544, -5.0220144e-05, -2.321794e-06, -2.7163756e-05, 0.00083960575, -5.850646e-05, -1.652374e-06, 0.00038475564, 0.0008068475, -6.618562e-05, -9.250065e-07, 0.0007784943, 0.0007669673, -7.316853e-05, -1.497222e-07, 0.0011506232, 0.00072050426, -7.937563e-05, 6.629815e-07, 0.0014979994, 0.000668063, -8.473774e-05, 1.5022744e-06, 0.0018177973, 0.0006103056, -8.919661e-05, 2.3571292e-06, 0.0021075346, 0.000547943, -9.270552e-05, 3.2164576e-06, 0.002365095, 0.00048172637, -9.522962e-05, 4.069244e-06, 0.002588746, 0.00041243774, -9.674611e-05, 4.9046766e-06, 0.0027771518, 0.00034088065, -9.7244396e-05, 5.7122747e-06, 0.0029293816, 0.00026787055, -9.672597e-05, 6.482007e-06, 0.0030449138, 0.00019422543, -9.520421e-05, 7.204406e-06, 0.0031236338, 0.00012075634, -9.270407e-05, 7.870673e-06, 0.0031658295, 4.8258335e-05, -8.926157e-05, 8.472772e-06, 0.0031721801, -2.2498389e-05, -8.492326e-05, 9.003513e-06, 0.003143742, -9.077683e-05, -7.974546e-05, 9.4566285e-06, 0.0030819303, -0.00015588106, -7.379349e-05, 9.826832e-06, 0.0029884963, -0.00021716346, -6.714076e-05, 1.0109866e-05, 0.0028655012, -0.00027403128, -5.9867805e-05, 1.030254e-05, 0.0027152882, -0.00032595254, -5.206122e-05, 1.0402753e-05, 0.0025404498, -0.000372461, -4.3812594e-05, 1.04095e-05, 0.0023437948, -0.0004131604, -3.5217337e-05, 1.032287e-05, 0.0021283112, -0.0004477277, -2.6373558e-05, 1.0144035e-05, 0.0018971302, -0.0004759157, -1.738085e-05, 9.875211e-06, 0.0016534871, -0.0004975543, -8.339134e-06, 9.5196265e-06, 0.001400683, -0.0005125514, 6.5249236e-07, 9.081469e-06, 0.0011420455, -0.00052089227, 9.4969e-06, 8.565822e-06, 0.00088089047, -0.00052263855, 1.810001e-05, 7.978593e-06, 0.00062048424, -0.0005179262, 2.6371838e-05, 7.3264337e-06, 0.00036400717, -0.0005069625, 3.422745e-05, 6.6166567e-06, 0.00011451893, -0.00049002253, 4.1587886e-05, 5.8571363e-06, -0.0001250745, -0.0004674449, 4.8380953e-05, 5.0562144e-06, -0.0003520511, -0.00043962628, 5.4541957e-05, 4.222595e-06, -0.0005639008, -0.00040701643, 6.0014332e-05, 3.365242e-06, -0.00075835024, -0.0003701115, 6.475016e-05, 2.4932692e-06, -0.0009333844, -0.00032944788, 6.871057e-05, 1.6158366e-06, -0.0010872651, -0.00028559507, 7.186606e-05, 7.4204394e-07, -0.0012185457, -0.00023914858, 7.419667e-05, -1.1917229e-07, -0.0013260824, -0.00019072261, 7.5692085e-05, -9.591386e-07, -0.0014090413, -0.00014094257, 7.635154e-05, -1.7695393e-06, -0.0014669029, -9.043767e-05, 7.6183744e-05, -2.5425059e-06, -0.0014994614, -3.9833558e-05, 7.5206575e-05, -3.2706998e-06, -0.0015068215, 1.0254878e-05, 7.344675e-05, -3.9473884e-06, -0.0014893912, 5.9230428e-05, 7.093935e-05, -4.566511e-06, -0.0014478713, 0.00010652019, 6.772732e-05, -5.122739e-06, -0.0013832418, 0.00015158176, 6.386082e-05, -5.6115227e-06, -0.0012967449, 0.00019390904, 5.93965e-05, -6.0291327e-06, -0.0011898658, 0.00023303744, 5.4396824e-05, -6.372689e-06, -0.0010643104, 0.00026854855, 4.8929178e-05, -6.6401776e-06, -0.0009219817, 0.0003000742, 4.3065043e-05, -6.830463e-06, -0.0007649533, 0.00032729987, 3.6879126e-05, -6.943284e-06, -0.00059544214, 0.00034996742, 3.0448418e-05, -6.9792427e-06, -0.00041577968, 0.00036787707, 2.3851286e-05, -6.9397847e-06, -0.0002283824, 0.00038088873, 1.716655e-05, -6.827166e-06, -3.5721743e-05, 0.0003889226, 1.0472569e-05, -6.6444177e-06, 0.00015970602, 0.00039195913, 3.84635e-06, -6.3952925e-06, 0.0003554097, 0.00039003804, -2.637314e-06, -6.0842167e-06, 0.0005489325, 0.000383257, -8.906665e-06, -5.7162215e-06, 0.0007378806, 0.00037176942, -1.4893752e-05, -5.2968808e-06, 0.00091995014, 0.0003557817, -2.0535148e-05, -4.8322336e-06, 0.0010929531, 0.00033554994, -2.5772597e-05, -4.328711e-06, 0.0012548412, 0.00031137612, -3.0553598e-05, -3.7930529e-06, 0.0014037276, 0.00028360382, -3.483191e-05, -3.2322278e-06, 0.0015379067, 0.00025261342, -3.8567974e-05, -2.653347e-06, 0.0016558714, 0.00021881713, -4.172925e-05, -2.0635835e-06, 0.0017563275, 0.00018265363, -4.4290467e-05, -1.4700853e-06, 0.0018382053, 0.0001445825, -4.6233796e-05, -8.798973e-07, 0.0019006693, 0.00010507852, -4.7548918e-05, -2.9988044e-07, 0.001943124, 6.462584e-05, -4.8233018e-05, 2.63363e-07, 0.0019652168, 2.3712253e-05, -4.829067e-05, 8.035608e-07, 0.001966839, -1.7176591e-05, -4.7733673e-05, 1.3148367e-06, 0.0019481225, -5.7562815e-05, -4.6580783e-05, 1.7917708e-06, 0.001909436, -9.6981734e-05, -4.4857356e-05, 2.229454e-06, 0.0018513753, -0.00013498706, -4.2594966e-05, 2.6235343e-06, 0.0017747541, -0.00017115581, -3.983091e-05, 2.9702587e-06, 0.0016805907, -0.00020509283, -3.6607682e-05, 3.2665032e-06, 0.0015700932, -0.00023643493, -3.2972388e-05, 3.5097996e-06, 0.0014446424, -0.00026485464, -2.8976121e-05, 3.6983504e-06, 0.0013057735, -0.00029006338, -2.4673294e-05, 3.8310386e-06, 0.0011551554, -0.0003118142, -2.012095e-05, 3.907428e-06, 0.0009945696, -0.00032990403, -1.537806e-05, 3.9277547e-06, 0.00082588807, -0.00034417518, -1.0504799e-05, 3.892914e-06, 0.0006510498, -0.0003545167, -5.5618216e-06, 3.8044357e-06, 0.00047203756, -0.0003608646, -6.095561e-07, 3.6644583e-06, 0.0002908543, -0.0003632021, 4.2925003e-06, 3.4756895e-06, 0.00010949978, -0.0003615589, 9.086454e-06, 3.2413664e-06, -7.005265e-05, -0.00035601013, 1.3716667e-05, 2.9652074e-06, -0.00024587815, -0.00034667485, 1.8130359e-05, 2.6513612e-06, -0.000416122, -0.00033371375, 2.2278178e-05, 2.3043497e-06, -0.00057901966, -0.00031732683, 2.6114716e-05, 1.929009e-06, -0.0007329159, -0.00029775038, 2.959897e-05, 1.5304275e-06, -0.00087628193, -0.00027525355, 3.269475e-05, 1.1138819e-06, -0.0010077311, -0.00025013494, 3.5371e-05, 6.847718e-07, -0.0011260324, -0.00022271842, 3.760211e-05, 2.4855487e-07, -0.0012301225, -0.00019334916, 3.936808e-05, -1.893183e-07, -0.001319115, -0.00016238925, 4.0654697e-05, -6.234677e-07, -0.0013923077, -0.0001302132, 4.1453575e-05, -1.0486458e-06, -0.0014491879, -9.720347e-05, 4.1762174e-05, -1.4597965e-06, -0.0014894352, -6.374589e-05, 4.1583724e-05, -1.8521115e-06, -0.0015129221, -3.0225176e-05, 4.092709e-05, -2.221082e-06, -0.0015197119, 2.9794865e-06, 3.980659e-05, -2.5625463e-06, -0.0015100557, 3.5498742e-05, 3.8241713e-05, -2.8727338e-06, -0.0014843857, 6.697716e-05, 3.6256835e-05, -3.1483007e-06, -0.0014433075, 9.707708e-05, 3.388084e-05, -3.386364e-06, -0.0013875904, 0.00012548224, 3.1146705e-05, -3.584526e-06, -0.0013181557, 0.00015190107, 2.8091063e-05, -3.740896e-06, -0.0012360639, 0.00017606962, 2.4753714e-05, -3.854103e-06, -0.0011424997, 0.00019775413, 2.1177106e-05, -3.9233023e-06, -0.0010387572, 0.00021675328, 1.74058e-05, -3.9481793e-06, -0.0009262218, 0.00023289995, 1.3485926e-05, -3.928943e-06, -0.0008063545, 0.00024606255, 9.464609e-06, -3.866315e-06, -0.0006806726, 0.00025614596, 5.3894196e-06, -3.7615139e-06, -0.0005507317, 0.00026309196, 1.3078055e-06, -3.6162312e-06, -0.00041810746, 0.00026687945, -2.7334515e-06, -3.4326067e-06, -0.00028437664, 0.00026752386, -6.688769e-06, -3.2131943e-06, -0.00015109948, 0.0002650765, -1.0514272e-05, -2.9609264e-06, -1.9801768e-05, 0.00025962334, -1.4168271e-05, -2.6790735e-06, 0.00010804198, 0.00025128332, -1.7611716e-05, -2.3712018e-06, 0.00023102465, 0.00024020665, -2.0808595e-05, -2.041126e-06, 0.0003478215, 0.00022657229, -2.3726312e-05, -1.6928611e-06, 0.000457204, 0.0002105856, -2.6336e-05, -1.3305736e-06, 0.00055805227, 0.0001924754, -2.86128e-05, -9.585298e-07, 0.0006493661, 0.00017249103, -3.053608e-05, -5.8104513e-07, 0.0007302744, 0.00015089898, -3.2089603e-05, -2.0243363e-07, 0.00080004294, 0.0001279797, -3.3261647e-05, 1.7304232e-07, 0.00085808046, 0.00010402399, -3.4045068e-05, 5.412203e-07, 0.000903943, 7.932951e-05, -3.4437293e-05, 8.9808447e-07, 0.0009373362, 5.4197226e-05, -3.4440294e-05, 1.2398096e-06, 0.00095811655, 2.8927887e-05, -3.4060486e-05, 1.5628023e-06, 0.00096629, 3.8185226e-06, -3.3308566e-05, 1.8637385e-06, 0.0009620094, -2.0840904e-05, -3.219934e-05, 2.139598e-06, 0.0009455702, -4.477073e-05, -3.075146e-05, 2.3876942e-06, 0.0009174042, -6.770467e-05, -2.8987177e-05, 2.6056998e-06, 0.00087807275, -8.939263e-05, -2.6931988e-05, 2.7916674e-06, 0.00082825747, -0.00010960339, -2.461432e-05, 2.9440466e-06, 0.0007687504, -0.00012812686, -2.2065136e-05, 3.0616948e-06, 0.0007004428, -0.00014477625, -1.9317536e-05, 3.1438838e-06, 0.0006243134, -0.00015938978, -1.6406348e-05, 3.1903023e-06, 0.000541415, -0.00017183211, -1.33676895e-05, 3.2010514e-06, 0.0004528613, -0.00018199554, -1.0238536e-05, 3.1766376e-06, 0.00035981278, -0.00018980069, -7.0562724e-06, 3.1179597e-06, 0.00026346243, -0.00019519699, -3.8582616e-06, 3.0262931e-06, 0.00016502131, -0.00019816274, -6.8140974e-07, 2.9032674e-06, 6.570411e-05, -0.00019870495, 2.4382505e-06, 2.7508431e-06, -3.3284992e-05, -0.00019685866, 5.465961e-06, 2.5712827e-06, -0.0001307662, -0.00019268612, 8.368619e-06, 2.3671205e-06, -0.00022559743, -0.0001862756, 1.111513e-05, 2.1411277e-06, -0.0003166869, -0.00017773996, 1.3676734e-05, 1.896278e-06, -0.00040300505, -0.00016721482, 1.6027298e-05, 1.635709e-06, -0.00048359542, -0.00015485672, 1.814357e-05, 1.3626835e-06, -0.0005575847, -0.00014084089, 2.0005407e-05, 1.0805502e-06, -0.00062419113, -0.00012535887, 2.1595948e-05, 7.927032e-07, -0.0006827326, -0.000108616085, 2.2901751e-05, 5.025426e-07, -0.0007326324, -9.082921e-05, 2.3912902e-05, 2.1343516e-07, -0.0007734245, -7.222342e-05, 2.4623056e-05, -7.132415e-08, -0.00080475706, -5.3029675e-05, 2.502946e-05, -3.4854867e-07, -0.0008263945, -3.3481938e-05, 2.513292e-05, -6.1519495e-07, -0.0008382184, -1.3814398e-05, 2.4937726e-05, -8.6839543e-07, -0.00084022695, 5.7412394e-06, 2.445156e-05, -1.1054885e-06, -0.000832533, 2.4958403e-05, 2.3685325e-05, -1.3240457e-06, -0.0008153609, 4.36182e-05, 2.2652985e-05, -1.5218957e-06, -0.00078904204, 6.151183e-05, 2.1371345e-05, -1.6971446e-06, -0.0007540092, 7.844284e-05, 1.98598e-05, -1.8481938e-06, -0.0007107897, 9.4229166e-05, 1.8140086e-05, -1.973753e-06, -0.0006599982, 0.00010870506, 1.6235963e-05, -2.072849e-06, -0.0006023276, 0.00012172271, 1.4172929e-05, -2.1448332e-06, -0.0005385399, 0.00013315363, 1.197788e-05, -2.189382e-06, -0.0004694564, 0.0001428899, 9.678783e-06, -2.2064958e-06, -0.00039594696, 0.000150845, 7.3043298e-06, -2.1964927e-06, -0.0003189192, 0.00015695447, 4.8835964e-06, -2.16e-06, -0.00023930735, 0.00016117636, 2.4456945e-06, -2.0979417e-06, -0.000158061, 0.00016349126, 1.9438557e-08, -2.0115217e-06, -7.613381e-05, 0.00016390221, -2.3669863e-06, -1.9022065e-06, 5.5276073e-06, 0.00016243423, -4.6863383e-06, -1.7717024e-06, 8.599451e-05, 0.00015913373, -6.91262e-06, -1.6219325e-06, 0.00016436652, 0.00015406757, -9.021357e-06, -1.4550101e-06, 0.0002397816, 0.000147322, -1.09898565e-05, -1.2732113e-06, 0.00031142536, 0.00013900126, -1.2797443e-05, -1.0789458e-06, 0.00037853981, 0.00012922616, -1.4425657e-05, -8.7472654e-07, 0.0004404311, 0.000118132346, -1.585844e-05, -6.631388e-07, 0.0004964765, 0.000105868516, -1.7082273e-05, -4.4680903e-07, 0.0005461306, 9.259446e-05, -1.8086295e-05, -2.2837375e-07, 0.0005889301, 7.847905e-05, -1.8862385e-05, -1.0448686e-08, 0.00062449806, 6.369811e-05, -1.94052e-05, 2.0440125e-07, 0.00065254676, 4.84323e-05, -1.9712208e-05, 4.1369077e-07, 0.0006728795, 3.2864893e-05, -1.9783653e-05, 6.150418e-07, 0.0006853914, 1.7179666e-05, -1.9622514e-05, 8.062092e-07, 0.00069006934, 1.5587267e-06, -1.9234425e-05, 9.851045e-07, 0.00068699016, -1.3819545e-05, -1.8627563e-05, 1.1498179e-06, 0.0006763186, -2.8782508e-05, -1.7812508e-05, 1.2986367e-06, 0.00065830396, -4.316516e-05, -1.6802087e-05, 1.4300626e-06, 0.0006332757, -5.6811925e-05, -1.5611182e-05, 1.5428252e-06, 0.0006016385, -6.957828e-05, -1.4256523e-05, 1.6358925e-06, 0.000563866, -8.1332255e-05, -1.2756469e-05, 1.7084797e-06, 0.00052049453, -9.195575e-05, -1.1130761e-05, 1.7600535e-06, 0.00047211576, -0.00010134568, -9.4002735e-06, 1.7903343e-06, 0.00041936894, -0.00010941489, -7.5867533e-06, 1.7992952e-06, 0.00036293277, -0.000116092924, -5.712553e-06, 1.7871583e-06, 0.00030351683, -0.00012132655, -3.8003616e-06, 1.7543875e-06, 0.00024185305, -0.00012508009, -1.8729359e-06, 1.7016795e-06, 0.00017868665, -0.00012733552, 4.716473e-08, 1.6299514e-06, 0.00011476754, -0.00012809242, 1.9378356e-06, 1.540327e-06, 5.0841467e-05, -0.0001273677, 3.7776758e-06, 1.43412e-06, -1.2358492e-05, -0.00012519505, 5.5462247e-06, 1.3128151e-06, -7.412017e-05, -0.000121624274, 7.224183e-06, 1.1780489e-06, -0.0001337602, -0.00011672055, 8.793616e-06, 1.0315878e-06, -0.00019063136, -0.00011056328, 1.0238141e-05, 8.753053e-07, -0.00024412952, -0.00010324503, 1.154309e-05, 7.1115886e-07, -0.00029369982, -9.487021e-05, 1.269565e-05, 5.4116543e-07, -0.00033884228, -8.555365e-05, 1.3684982e-05, 3.673775e-07, -0.00037911665, -7.541913e-05, 1.4502314e-05, 1.918583e-07, -0.00041414646, -6.459776e-05, 1.5141006e-05, 1.6657985e-08, -0.00044362227, -5.322641e-05, 1.5596595e-05, -1.5621004e-07, -0.00046730423, -4.1445935e-05, 1.5866808e-05, -3.2479178e-07, -0.00048502345, -2.9399558e-05, 1.5951551e-05, -4.872143e-07, -0.000496683, -1.7231143e-05, 1.5852878e-05, -6.417063e-07, -0.00050225767, -5.0835165e-06, 1.5574926e-05, -7.866165e-07, -0.000501793, 6.9031535e-06, 1.5123837e-05, -9.204313e-07, -0.00049540366, 1.8592944e-05, 1.4507653e-05, -1.0417896e-06, -0.00048327097, 2.985567e-05, 1.37361885e-05, -1.1494964e-06, -0.00046563946, 4.0568302e-05, 1.2820891e-05, -1.2425335e-06, -0.00044281324, 5.061626e-05, 1.17746795e-05, -1.3200689e-06, -0.00041515133, 5.989461e-05, 1.0611769e-05, -1.3814628e-06, -0.00038306252, 6.830909e-05, 9.347489e-06, -1.4262722e-06, -0.00034699994, 7.5777054e-05, 7.998085e-06, -1.4542526e-06, -0.00030745493, 8.22282e-05, 6.580511e-06, -1.4653576e-06, -0.0002649508, 8.760522e-05, 5.1122324e-06, -1.4597363e-06, -0.00022003613, 9.186418e-05, 3.6110046e-06, -1.437728e-06, -0.00017327811, 9.4974865e-05, 2.0946684e-06, -1.3998554e-06, -0.00012525555, 9.692086e-05, 5.8094145e-07, -1.3468156e-06, -7.655202e-05, 9.769953e-05, -9.127852e-07, -1.2794687e-06, -2.7749007e-05, 9.732179e-05, -2.3696427e-06, -1.198826e-06, 2.058078e-05, 9.581178e-05, -3.7734703e-06, -1.1060347e-06, 6.7879904e-05, 9.320637e-05, -5.1089905e-06, -1.0023633e-06, 0.000113612405, 8.955446e-05, -6.3619723e-06, -8.8918443e-07, 0.00015726963, 8.491628e-05, -7.5193757e-06, -7.6795754e-07, 0.00019837571, 7.9362464e-05, -8.569485e-06, -6.402103e-07, 0.00023649246, 7.2973075e-05, -9.502019e-06, -5.075201e-07, 0.00027122386, 6.5836495e-05, -1.0308231e-05, -3.7149482e-07, 0.00030221997, 5.8048292e-05, -1.0980981e-05, -2.3375374e-07, 0.0003291801, 4.970997e-05, -1.1514789e-05, -9.590874e-08, 0.0003518556, 4.09277e-05, -1.1905875e-05, 4.045425e-08, 0.0003700517, 3.1811025e-05, -1.2152172e-05, 1.7379317e-07, 0.0003836291, 2.247151e-05, -1.2253321e-05, 3.026269e-07, 0.00039250444, 1.3021434e-05, -1.2210649e-05, 4.2555126e-07, 0.00039665043, 3.5724718e-06, -1.2027122e-05, 5.4125417e-07, 0.00039609513, -5.7655866e-06, -1.1707282e-05, 6.48529e-07, 0.00039092085, -1.488608e-05, -1.1257177e-05, 7.46287e-07, 0.00038126216, -2.3686656e-05, -1.06842535e-05, 8.3356764e-07, 0.00036730347, -3.2070388e-05, -9.997255e-06, 9.095478e-07, 0.00034927618, -3.99468e-05, -9.206096e-06, 9.735488e-07, 0.00032745497, -4.7232814e-05, -8.32173e-06, 1.0250419e-06, 0.00030215413, -5.3853582e-05, -7.3560022e-06, 1.0636519e-06, 0.00027372318, -5.9743223e-05, -6.3214984e-06, 1.0891589e-06, 0.00024254216, -6.484542e-05, -5.231389e-06, 1.1014981e-06, 0.00020901674, -6.911395e-05, -4.0992645e-06, 1.1007583e-06, 0.00017357318, -7.2512994e-05, -2.9389716e-06, 1.0871773e-06, 0.00013665296, -7.501741e-05, -1.7644494e-06, 1.0611384e-06, 9.87074e-05, -7.6612865e-05, -5.895656e-07, 1.0231615e-06, 6.0192346e-05, -7.729579e-05, 5.720419e-07, 9.738964e-07, 2.1562724e-05, -7.707322e-05, 1.70712e-06, 9.141121e-07, -1.6732654e-05, -7.596262e-05, 2.802946e-06, 8.446863e-07, -5.425622e-05, -7.399141e-05, 3.8474677e-06, 7.6659353e-07, -9.058652e-05, -7.119654e-05, 4.82943e-06, 6.808917e-07, -0.00012532285, -6.762388e-05, 5.7384927e-06, 5.887091e-07, -0.0001580895, -6.332756e-05, 6.565335e-06, 4.912297e-07, -0.00018853977, -5.8369184e-05, 7.3017445e-06, 3.8967877e-07, -0.00021635942, -5.2817e-05, 7.940697e-06, 2.8530778e-07, -0.00024126982, -4.6744997e-05, 8.476415e-06, 1.7937968e-07, -0.00026303058, -4.0231964e-05, 8.904414e-06, 7.3153934e-08, -0.00028144172, -3.3360477e-05, 9.221534e-06, -3.2127932e-08, -0.00029634527, -2.6215896e-05, 9.425953e-06, -1.3525641e-07, -0.00030762635, -1.8885325e-05, 9.517186e-06, -2.350675e-07, -0.00031521395, -1.1456575e-05, 9.496067e-06, -3.3045538e-07, -0.0003190809, -4.017131e-06, 9.3647195e-06, -4.2038428e-07, -0.00031924344, 3.3468475e-06, 9.126507e-06, -5.038993e-07, -0.00031576038, 1.0551507e-05, 8.785978e-06, -5.80136e-07, -0.00030873172, 1.7516233e-05, 8.348788e-06, -6.48329e-07, -0.00029829674, 2.4164523e-05, 7.821619e-06, -7.0781925e-07, -0.00028463174, 3.042481e-05, 7.2120833e-06, -7.580597e-07, -0.00026794747, 3.6231206e-05, 6.5286226e-06, -7.9861974e-07, -0.00024848603, 4.152417e-05, 5.7803913e-06, -8.291885e-07, -0.0002265176, 4.625109e-05, 4.9771434e-06, -8.4957605e-07, -0.0002023368, 5.036678e-05, 4.1291064e-06, -8.597141e-07, -0.00017625892, 5.383387e-05, 3.2468565e-06, -8.59654e-07, -0.00014861595, 5.6623125e-05, 2.3411897e-06, -8.4956497e-07, -0.00011975233, 5.8713624e-05, 1.4229928e-06, -8.2972946e-07, -9.002095e-05, 6.0092883e-05, 5.031167e-07, -8.005384e-07, -5.977878e-05, 6.0756858e-05, -4.0774938e-07, -7.624847e-07, -2.9382736e-05, 6.0709834e-05, -1.2991989e-06, -7.161559e-07, 8.14462e-07, 5.9964248e-05, -2.1612236e-06, -6.622257e-07, 3.0468289e-05, 5.8540416e-05, -2.9843227e-06, -6.0144475e-07, 5.9246275e-05, 5.6466146e-05, -3.7596046e-06, -5.346306e-07, 8.6831635e-05, 5.377632e-05, -4.4788794e-06, -4.6265728e-07, 0.000112926675, 5.0512335e-05, -5.1347433e-06, -3.86444e-07, 0.00013725593, 4.6721547e-05, -5.7206485e-06, -3.0694392e-07, 0.00015956897, 4.2456617e-05, -6.230967e-06, -2.2513252e-07, 0.00017964284, 3.777479e-05, -6.6610396e-06, -1.4199584e-07, 0.00019728423, 3.2737193e-05, -7.0072147e-06, -5.8518935e-08, 0.0002123312, 2.7408027e-05, -7.2668718e-06, 2.4325521e-08, 0.00022465452, 2.1853803e-05, -7.438435e-06, 1.0558829e-07, 0.00023415861, 1.6142507e-05, -7.5213766e-06, 1.8435419e-07, 0.00024078209, 1.0342813e-05, -7.516201e-06, 2.597521e-07, 0.0002444979, 4.523257e-06, -7.4244263e-06, 3.3096438e-07, 0.0002453131, -1.2485418e-06, -7.2485464e-06, 3.9723534e-07, 0.00024326815, -6.9066514e-06, -6.991987e-06, 4.5787905e-07, 0.00023843585, -1.2387563e-05, -6.6590515e-06, 5.1228614e-07, 0.00023092006, -1.7630884e-05, -6.2548543e-06, 5.599294e-07, 0.0002208539, -2.2579985e-05, -5.7852503e-06, 6.0036876e-07, 0.00020839775, -2.718259e-05, -5.256753e-06, 6.3325484e-07, 0.0001937369, -3.139131e-05, -4.676449e-06, 6.583313e-07, 0.00017707904, -3.516412e-05, -4.051906e-06, 6.754366e-07, 0.00015865147, -3.846473e-05, -3.3910783e-06, 6.84504e-07, 0.00013869806, -4.1262923e-05, -2.702206e-06, 6.8556096e-07, 0.00011747629, -4.3534823e-05, -1.9937172e-06, 6.78727e-07, 9.5253905e-05, -4.526303e-05, -1.274126e-06, 6.642111e-07, 7.2305746e-05, -4.6436733e-05, -5.5193306e-07, 6.423075e-07, 4.891038e-05, -4.705172e-05, 1.6447315e-07, 6.133911e-07, 2.5346864e-05, -4.7110312e-05, 8.6691074e-07, 5.779116e-07, 1.8914722e-06, -4.662124e-05, 1.5474963e-06, 5.363872e-07, -2.1185442e-05, -4.559942e-05, 2.1987307e-06, 4.893973e-07, -4.3622476e-05, -4.4065688e-05, 2.81358e-06, 4.375749e-07, -6.517005e-05, -4.204645e-05, 3.3855483e-06, 3.815984e-07, -8.55931e-05, -3.9573297e-05, 3.9087445e-06, 3.2218284e-07, -0.00010467357, -3.668254e-05, 4.37794e-06, 2.6007118e-07, -0.00012221262, -3.341471e-05, 4.788619e-06, 1.9602507e-07, -0.00013803263, -2.9814035e-05, 5.137018e-06, 1.3081595e-07, -0.00015197888, -2.5927835e-05, 5.420156e-06, 6.521575e-08, -0.000163921, -2.1805956e-05, 5.6358576e-06, -1.1952672e-11, -0.000173754, -1.7500131e-05, 5.7827638e-06, -6.4120634e-08, -0.00018139913, -1.3063353e-05, 5.860334e-06, -1.263892e-07, -0.0001868043, -8.549245e-06, 5.8688393e-06, -1.8612985e-07, -0.00018994427, -4.011421e-06, 5.8093447e-06, -2.4269556e-07, -0.00019082046, 4.971275e-07, 5.683684e-06, -2.9548684e-07, -0.00018946052, 4.924638e-06, 5.494426e-06, -3.4395785e-07, -0.00018591754, 9.221154e-06, 5.2448327e-06, -3.8762184e-07, -0.00018026902, 1.3339076e-05, 4.9388077e-06, -4.2605583e-07, -0.0001726156, 1.7233668e-05, 4.580844e-06, -4.589044e-07, -0.00016307941, 2.0863534e-05, 4.1759586e-06, -4.8588265e-07, -0.00015180242, 2.4191033e-05, 3.7296281e-06, -5.0677835e-07, -0.00013894434, 2.7182663e-05, 3.2477167e-06, -5.214532e-07, -0.00012468056, 2.9809366e-05, 2.7364015e-06, -5.2984313e-07, -0.00010919985, 3.2046803e-05, 2.202096e-06, -5.319579e-07, -9.27019e-05, 3.3875545e-05, 1.651373e-06, -5.278795e-07, -7.5394855e-05, 3.5281228e-05, 1.090884e-06, -5.177603e-07, -5.7492776e-05, 3.625462e-05, 5.272819e-07, -5.018201e-07, -3.921303e-05, 3.679166e-05, -3.285569e-08, -4.803421e-07, -2.0773752e-05, 3.6893394e-05, -5.83102e-07, -4.5366892e-07, -2.3912733e-06, 3.6565907e-05, -1.1172526e-06, -4.221975e-07, 1.5722333e-05, 3.5820143e-05, -1.6293935e-06, -3.8637359e-07, 3.336164e-05, 3.4671713e-05, -2.113965e-06, -3.466858e-07, 5.033014e-05, 3.3140623e-05, -2.5658196e-06, -3.0365925e-07, 6.644237e-05, 3.1250976e-05, -2.9802754e-06, -2.5784885e-07, 8.152586e-05, 2.9030636e-05, -3.3531614e-06, -2.0983232e-07, 9.542295e-05, 2.6510814e-05, -3.6808583e-06, -1.6020327e-07, 0.00010799231, 2.3725677e-05, -3.960331e-06, -1.0956389e-07, 0.00011911037, 2.0711894e-05, -4.189153e-06, -5.8517998e-08, 0.0001286724, 1.750816e-05, -4.365525e-06, -7.663899e-09, 0.00013659344, 1.41547325e-05, -4.488286e-06, 4.2412374e-08, 0.00014280893, 1.0692924e-05, -4.556914e-06, 9.114367e-08, 0.00014727515, 7.1646145e-06, -4.5715233e-06, 1.3798794e-07, 0.00014996933, 3.6117533e-06, -4.5328516e-06, 1.8243412e-07, 0.00015088962, 7.587294e-08, -4.4422413e-06, 2.2400754e-07, 0.00015005471, -3.4023838e-06, -4.301613e-06, 2.622747e-07, 0.0001475033, -6.7837195e-06, -4.1134344e-06, 2.968478e-07, 0.00014329332, -1.0030616e-05, -3.880684e-06, 3.2738822e-07, 0.00013750092, -1.3107738e-05, -3.6068036e-06, 3.536098e-07, 0.00013021928, -1.5982303e-05, -3.2956561e-06, 3.752812e-07, 0.00012155731, -1.8624423e-05, -2.9514704e-06, 3.9222766e-07, 0.00011163802, -2.1007401e-05, -2.5787865e-06, 4.043321e-07, 0.00010059696, -2.3107985e-05, -2.182399e-06, 4.1153544e-07, 8.8580375e-05, -2.4906572e-05, -1.7672962e-06, 4.138364e-07, 7.574336e-05, -2.6387395e-05, -1.3386002e-06, 4.1129053e-07, 6.2247935e-05, -2.7538621e-05, -9.0150434e-07, 4.0400852e-07, 4.826102e-05, -2.8352426e-05, -4.6121215e-07, 3.9215408e-07, 3.395243e-05, -2.8825028e-05, -2.2877371e-08, 3.759412e-07, 1.9492882e-05, -2.8956656e-05, 4.0845538e-07, 3.5563068e-07, 5.0519816e-06, -2.8751478e-05, 8.279069e-07, 3.315265e-07, -9.203712e-06, -2.8217493e-05, 1.2308172e-06, 3.0397143e-07, -2.3112565e-05, -2.7366372e-05, 1.6127958e-06, 2.7334247e-07, -3.6519654e-05, -2.6213258e-05, 1.9697682e-06, 2.4004595e-07, -4.9278453e-05, -2.4776538e-05, 2.298017e-06, 2.045123e-07, -6.125238e-05, -2.3077575e-05, 2.5942204e-06, 1.6719062e-07, -7.2316216e-05, -2.1140404e-05, 2.8554823e-06, 1.2854323e-07, -8.2357365e-05, -1.8991419e-05, 3.0793606e-06, 8.904007e-08, -9.127695e-05, -1.6659023e-05, 3.2638857e-06, 4.9153147e-08, -9.899071e-05, -1.4173269e-05, 3.4075777e-06, 9.350997e-09, -0.00010542977, -1.1565476e-05, 3.509453e-06, -2.9906634e-08, -0.000110541114, -8.8678535e-06, 3.5690296e-06, -6.8173996e-08, -0.000114288, -6.113115e-06, 3.5863227e-06, -1.05024256e-07, -0.00011665008, -3.3340827e-06, 3.561837e-06, -1.4005413e-07, -0.00011762337, -5.6331345e-07, 3.4965524e-06, -1.7288812e-07, -0.000117220006, 2.1672777e-06, 3.3919043e-06, -2.0318245e-07};
	localparam real hb[0:1999] = {0.024986578, 0.000116877105, -3.896343e-05, -2.2712003e-07, 0.024869869, 0.0003495672, -3.6725352e-05, -6.683011e-07, 0.02463752, 0.00057908345, -3.2282736e-05, -1.071189e-06, 0.02429164, 0.00080335606, -2.5699466e-05, -1.4122909e-06, 0.023835355, 0.0010203768, -1.7068134e-05, -1.6701244e-06, 0.023272775, 0.0012282217, -6.508329e-06, -1.825436e-06, 0.02260895, 0.0014250721, 5.835373e-06, -1.8613864e-06, 0.021849804, 0.0016092348, 1.979567e-05, -1.7637041e-06, 0.021002075, 0.0017791594, 3.5185032e-05, -1.5208042e-06, 0.020073237, 0.0019334549, 5.1798383e-05, -1.1238726e-06, 0.019071415, 0.0020709035, 6.941594e-05, -5.669145e-07, 0.018005302, 0.0021904726, 8.7806206e-05, 1.5323168e-07, 0.016884053, 0.0022913238, 0.000106729, 1.0369153e-06, 0.015717195, 0.0023728213, 0.00012593858, 2.0817276e-06, 0.014514523, 0.0024345345, 0.00014518676, 3.2825897e-06, 0.01328599, 0.0024762424, 0.000164226, 4.6318687e-06, 0.012041612, 0.0024979326, 0.00018281244, 6.119525e-06, 0.010791358, 0.0024997983, 0.00020070883, 7.733287e-06, 0.009545049, 0.0024822343, 0.00021768737, 9.458844e-06, 0.008312262, 0.0024458296, 0.00023353235, 1.1280068e-05, 0.0071022296, 0.0023913574, 0.00024804258, 1.31792485e-05, 0.0059237573, 0.0023197657, 0.0002610337, 1.5137347e-05, 0.004785133, 0.0022321627, 0.00027234023, 1.7134254e-05, 0.003694055, 0.002129803, 0.00028181716, 1.9149073e-05, 0.0026575602, 0.0020140712, 0.0002893417, 2.116038e-05, 0.0016819648, 0.0018864649, 0.00029481426, 2.3146522e-05, 0.0007728115, 0.0017485761, 0.00029815955, 2.5085883e-05, -6.517271e-05, 0.0016020724, 0.00029932705, 2.6957157e-05, -0.0008281093, 0.0014486772, 0.0002982914, 2.8739623e-05, -0.0015129913, 0.0012901495, 0.00029505236, 3.0413386e-05, -0.002117696, 0.0011282647, 0.0002896347, 3.195963e-05, -0.0026409882, 0.00096479343, 0.0002820874, 3.3360822e-05, -0.003082513, 0.00080148317, 0.00027248287, 3.4600955e-05, -0.0034427792, 0.00064003846, 0.000260916, 3.5665686e-05, -0.0037231334, 0.0004821034, 0.00024750258, 3.6542533e-05, -0.003925726, 0.00032924407, 0.00023237792, 3.7221005e-05, -0.004053466, 0.00018293266, 0.00021569492, 3.76927e-05, -0.0041099745, 4.453296e-05, 0.00019762217, 3.79514e-05, -0.0040995227, -8.471297e-05, 0.00017834186, 3.7993144e-05, -0.0040269704, -0.00020369625, 0.00015804752, 3.7816237e-05, -0.0038976963, -0.00031145103, 0.00013694167, 3.742127e-05, -0.0037175252, -0.00040716256, 0.00011523339, 3.6811085e-05, -0.0034926496, -0.0004901733, 9.3135954e-05, 3.599074e-05, -0.0032295508, -0.00055998715, 7.086427e-05, 3.4967423e-05, -0.002934917, -0.0006162719, 4.8632493e-05, 3.3750366e-05, -0.0026155617, -0.0006588598, 2.6651622e-05, 3.235072e-05, -0.0022783414, -0.0006877456, 5.1271536e-06, 3.0781408e-05, -0.0019300748, -0.00070308376, -1.5743133e-05, 2.9056979e-05, -0.0015774649, -0.0007051833, -3.577129e-05, 2.7193415e-05, -0.0012270228, -0.00069450086, -5.4781158e-05, 2.5207955e-05, -0.00088499615, -0.00067163265, -7.261017e-05, 2.311889e-05, -0.00055730145, -0.0006373044, -8.911096e-05, 2.0945343e-05, -0.0002494623, -0.00059236056, -0.00010415277, 1.8707058e-05, 3.3447053e-05, -0.00053775206, -0.00011762269, 1.6424181e-05, 0.00028685166, -0.00047452268, -0.00012942658, 1.4117025e-05, 0.0005067189, -0.00040379557, -0.0001394899, 1.1805854e-05, 0.00068959437, -0.00032675808, -0.00014775814, 9.510665e-06, 0.0008326304, -0.00024464677, -0.00015419716, 7.2509692e-06, 0.0009336064, -0.00015873181, -0.00015879319, 5.0455933e-06, 0.0009909424, -7.03015e-05, -0.0001615527, 2.9124817e-06, 0.0010037036, 1.9353303e-05, -0.00016250192, 8.6851696e-07, 0.000971598, 0.00010895448, -0.00016168621, -1.0706473e-06, 0.00089496677, 0.00019725144, -0.00015916926, -2.890736e-06, 0.0007747661, 0.0002830354, -0.00015503199, -4.578985e-06, 0.0006125435, 0.0003651528, -0.0001493714, -6.1242554e-06, 0.00041040673, 0.00044251818, -0.00014229909, -7.517124e-06, 0.00017098685, 0.0005141254, -0.00013393987, -8.749958e-06, -0.000102604055, 0.0005790583, -0.00012442996, -9.816967e-06, -0.00040682033, 0.00063650013, -0.00011391535, -1.0714228e-05, -0.0007377343, 0.00068574096, -0.000102549915, -1.1439698e-05, -0.0010910918, 0.00072618475, -9.049353e-05, -1.1993197e-05, -0.0014623696, 0.0007573539, -7.791015e-05, -1.237638e-05, -0.0018468365, 0.0007788933, -6.496585e-05, -1.2592673e-05, -0.002239615, 0.0007905721, -5.1826923e-05, -1.2647208e-05, -0.0026357428, 0.0007922844, -3.8657945e-05, -1.2546729e-05, -0.0030302363, 0.00078404846, -2.5619947e-05, -1.22994825e-05, -0.0034181513, 0.0007660045, -1.2868641e-05, -1.1915097e-05, -0.0037946438, 0.0007384107, -5.527264e-07, -1.1404446e-05, -0.0041550267, 0.00070163846, 1.1187671e-05, -1.0779499e-05, -0.0044948263, 0.000656166, 2.2222448e-05, -1.0053163e-05, -0.004809833, 0.00060257106, 3.2432832e-05, -9.239121e-06, -0.005096149, 0.0005415224, 4.1712527e-05, -8.351654e-06, -0.0053502326, 0.00047377063, 4.9968694e-05, -7.4054738e-06, -0.0055689337, 0.0004001377, 5.7122783e-05, -6.415538e-06, -0.005749531, 0.00032150644, 6.311115e-05, -5.3968797e-06, -0.005889757, 0.00023880896, 6.788551e-05, -4.3644327e-06, -0.005987819, 0.00015301503, 7.1413204e-05, -3.33286e-06, -0.0060424167, 6.5120075e-05, 7.367729e-05, -2.3163923e-06, -0.0060527516, -2.3866987e-05, 7.467643e-05, -1.3286729e-06, -0.006018531, -0.00011293571, 7.442458e-05, -3.8261123e-07, -0.0059399647, -0.00020108608, 7.295059e-05, 5.097503e-07, -0.005817757, -0.00028734, 7.029756e-05, 1.3373586e-06, -0.0056530945, -0.00037075247, 6.652203e-05, 2.0902578e-06, -0.005447625, -0.00045042214, 6.169313e-05, 2.759682e-06, -0.0052034347, -0.00052550115, 5.589148e-05, 3.3381343e-06, -0.004923017, -0.00059520424, 4.9208058e-05, 3.819447e-06, -0.004609243, -0.00065881707, 4.1742933e-05, 4.198827e-06, -0.0042653196, -0.0007157032, 3.3603916e-05, 4.472884e-06, -0.003894752, -0.0007653107, 2.4905143e-05, 4.639643e-06, -0.0035012984, -0.0008071772, 1.5765636e-05, 4.698537e-06, -0.003088926, -0.0008409337, 6.307793e-06, 4.6503856e-06, -0.0026617618, -0.0008663077, -3.3441117e-06, 4.4973604e-06, -0.0022240446, -0.00088312494, -1.3065424e-05, 4.2429283e-06, -0.0017800763, -0.0008913099, -2.2732595e-05, 3.8917874e-06, -0.0013341709, -0.000890885, -3.2224616e-05, 3.4497868e-06, -0.0008906079, -0.00088196935, -4.142441e-05, 2.9238345e-06, -0.0004535831, -0.00086477544, -5.0220144e-05, 2.321794e-06, -2.7163756e-05, -0.00083960575, -5.850646e-05, 1.652374e-06, 0.00038475564, -0.0008068475, -6.618562e-05, 9.250065e-07, 0.0007784943, -0.0007669673, -7.316853e-05, 1.497222e-07, 0.0011506232, -0.00072050426, -7.937563e-05, -6.629815e-07, 0.0014979994, -0.000668063, -8.473774e-05, -1.5022744e-06, 0.0018177973, -0.0006103056, -8.919661e-05, -2.3571292e-06, 0.0021075346, -0.000547943, -9.270552e-05, -3.2164576e-06, 0.002365095, -0.00048172637, -9.522962e-05, -4.069244e-06, 0.002588746, -0.00041243774, -9.674611e-05, -4.9046766e-06, 0.0027771518, -0.00034088065, -9.7244396e-05, -5.7122747e-06, 0.0029293816, -0.00026787055, -9.672597e-05, -6.482007e-06, 0.0030449138, -0.00019422543, -9.520421e-05, -7.204406e-06, 0.0031236338, -0.00012075634, -9.270407e-05, -7.870673e-06, 0.0031658295, -4.8258335e-05, -8.926157e-05, -8.472772e-06, 0.0031721801, 2.2498389e-05, -8.492326e-05, -9.003513e-06, 0.003143742, 9.077683e-05, -7.974546e-05, -9.4566285e-06, 0.0030819303, 0.00015588106, -7.379349e-05, -9.826832e-06, 0.0029884963, 0.00021716346, -6.714076e-05, -1.0109866e-05, 0.0028655012, 0.00027403128, -5.9867805e-05, -1.030254e-05, 0.0027152882, 0.00032595254, -5.206122e-05, -1.0402753e-05, 0.0025404498, 0.000372461, -4.3812594e-05, -1.04095e-05, 0.0023437948, 0.0004131604, -3.5217337e-05, -1.032287e-05, 0.0021283112, 0.0004477277, -2.6373558e-05, -1.0144035e-05, 0.0018971302, 0.0004759157, -1.738085e-05, -9.875211e-06, 0.0016534871, 0.0004975543, -8.339134e-06, -9.5196265e-06, 0.001400683, 0.0005125514, 6.5249236e-07, -9.081469e-06, 0.0011420455, 0.00052089227, 9.4969e-06, -8.565822e-06, 0.00088089047, 0.00052263855, 1.810001e-05, -7.978593e-06, 0.00062048424, 0.0005179262, 2.6371838e-05, -7.3264337e-06, 0.00036400717, 0.0005069625, 3.422745e-05, -6.6166567e-06, 0.00011451893, 0.00049002253, 4.1587886e-05, -5.8571363e-06, -0.0001250745, 0.0004674449, 4.8380953e-05, -5.0562144e-06, -0.0003520511, 0.00043962628, 5.4541957e-05, -4.222595e-06, -0.0005639008, 0.00040701643, 6.0014332e-05, -3.365242e-06, -0.00075835024, 0.0003701115, 6.475016e-05, -2.4932692e-06, -0.0009333844, 0.00032944788, 6.871057e-05, -1.6158366e-06, -0.0010872651, 0.00028559507, 7.186606e-05, -7.4204394e-07, -0.0012185457, 0.00023914858, 7.419667e-05, 1.1917229e-07, -0.0013260824, 0.00019072261, 7.5692085e-05, 9.591386e-07, -0.0014090413, 0.00014094257, 7.635154e-05, 1.7695393e-06, -0.0014669029, 9.043767e-05, 7.6183744e-05, 2.5425059e-06, -0.0014994614, 3.9833558e-05, 7.5206575e-05, 3.2706998e-06, -0.0015068215, -1.0254878e-05, 7.344675e-05, 3.9473884e-06, -0.0014893912, -5.9230428e-05, 7.093935e-05, 4.566511e-06, -0.0014478713, -0.00010652019, 6.772732e-05, 5.122739e-06, -0.0013832418, -0.00015158176, 6.386082e-05, 5.6115227e-06, -0.0012967449, -0.00019390904, 5.93965e-05, 6.0291327e-06, -0.0011898658, -0.00023303744, 5.4396824e-05, 6.372689e-06, -0.0010643104, -0.00026854855, 4.8929178e-05, 6.6401776e-06, -0.0009219817, -0.0003000742, 4.3065043e-05, 6.830463e-06, -0.0007649533, -0.00032729987, 3.6879126e-05, 6.943284e-06, -0.00059544214, -0.00034996742, 3.0448418e-05, 6.9792427e-06, -0.00041577968, -0.00036787707, 2.3851286e-05, 6.9397847e-06, -0.0002283824, -0.00038088873, 1.716655e-05, 6.827166e-06, -3.5721743e-05, -0.0003889226, 1.0472569e-05, 6.6444177e-06, 0.00015970602, -0.00039195913, 3.84635e-06, 6.3952925e-06, 0.0003554097, -0.00039003804, -2.637314e-06, 6.0842167e-06, 0.0005489325, -0.000383257, -8.906665e-06, 5.7162215e-06, 0.0007378806, -0.00037176942, -1.4893752e-05, 5.2968808e-06, 0.00091995014, -0.0003557817, -2.0535148e-05, 4.8322336e-06, 0.0010929531, -0.00033554994, -2.5772597e-05, 4.328711e-06, 0.0012548412, -0.00031137612, -3.0553598e-05, 3.7930529e-06, 0.0014037276, -0.00028360382, -3.483191e-05, 3.2322278e-06, 0.0015379067, -0.00025261342, -3.8567974e-05, 2.653347e-06, 0.0016558714, -0.00021881713, -4.172925e-05, 2.0635835e-06, 0.0017563275, -0.00018265363, -4.4290467e-05, 1.4700853e-06, 0.0018382053, -0.0001445825, -4.6233796e-05, 8.798973e-07, 0.0019006693, -0.00010507852, -4.7548918e-05, 2.9988044e-07, 0.001943124, -6.462584e-05, -4.8233018e-05, -2.63363e-07, 0.0019652168, -2.3712253e-05, -4.829067e-05, -8.035608e-07, 0.001966839, 1.7176591e-05, -4.7733673e-05, -1.3148367e-06, 0.0019481225, 5.7562815e-05, -4.6580783e-05, -1.7917708e-06, 0.001909436, 9.6981734e-05, -4.4857356e-05, -2.229454e-06, 0.0018513753, 0.00013498706, -4.2594966e-05, -2.6235343e-06, 0.0017747541, 0.00017115581, -3.983091e-05, -2.9702587e-06, 0.0016805907, 0.00020509283, -3.6607682e-05, -3.2665032e-06, 0.0015700932, 0.00023643493, -3.2972388e-05, -3.5097996e-06, 0.0014446424, 0.00026485464, -2.8976121e-05, -3.6983504e-06, 0.0013057735, 0.00029006338, -2.4673294e-05, -3.8310386e-06, 0.0011551554, 0.0003118142, -2.012095e-05, -3.907428e-06, 0.0009945696, 0.00032990403, -1.537806e-05, -3.9277547e-06, 0.00082588807, 0.00034417518, -1.0504799e-05, -3.892914e-06, 0.0006510498, 0.0003545167, -5.5618216e-06, -3.8044357e-06, 0.00047203756, 0.0003608646, -6.095561e-07, -3.6644583e-06, 0.0002908543, 0.0003632021, 4.2925003e-06, -3.4756895e-06, 0.00010949978, 0.0003615589, 9.086454e-06, -3.2413664e-06, -7.005265e-05, 0.00035601013, 1.3716667e-05, -2.9652074e-06, -0.00024587815, 0.00034667485, 1.8130359e-05, -2.6513612e-06, -0.000416122, 0.00033371375, 2.2278178e-05, -2.3043497e-06, -0.00057901966, 0.00031732683, 2.6114716e-05, -1.929009e-06, -0.0007329159, 0.00029775038, 2.959897e-05, -1.5304275e-06, -0.00087628193, 0.00027525355, 3.269475e-05, -1.1138819e-06, -0.0010077311, 0.00025013494, 3.5371e-05, -6.847718e-07, -0.0011260324, 0.00022271842, 3.760211e-05, -2.4855487e-07, -0.0012301225, 0.00019334916, 3.936808e-05, 1.893183e-07, -0.001319115, 0.00016238925, 4.0654697e-05, 6.234677e-07, -0.0013923077, 0.0001302132, 4.1453575e-05, 1.0486458e-06, -0.0014491879, 9.720347e-05, 4.1762174e-05, 1.4597965e-06, -0.0014894352, 6.374589e-05, 4.1583724e-05, 1.8521115e-06, -0.0015129221, 3.0225176e-05, 4.092709e-05, 2.221082e-06, -0.0015197119, -2.9794865e-06, 3.980659e-05, 2.5625463e-06, -0.0015100557, -3.5498742e-05, 3.8241713e-05, 2.8727338e-06, -0.0014843857, -6.697716e-05, 3.6256835e-05, 3.1483007e-06, -0.0014433075, -9.707708e-05, 3.388084e-05, 3.386364e-06, -0.0013875904, -0.00012548224, 3.1146705e-05, 3.584526e-06, -0.0013181557, -0.00015190107, 2.8091063e-05, 3.740896e-06, -0.0012360639, -0.00017606962, 2.4753714e-05, 3.854103e-06, -0.0011424997, -0.00019775413, 2.1177106e-05, 3.9233023e-06, -0.0010387572, -0.00021675328, 1.74058e-05, 3.9481793e-06, -0.0009262218, -0.00023289995, 1.3485926e-05, 3.928943e-06, -0.0008063545, -0.00024606255, 9.464609e-06, 3.866315e-06, -0.0006806726, -0.00025614596, 5.3894196e-06, 3.7615139e-06, -0.0005507317, -0.00026309196, 1.3078055e-06, 3.6162312e-06, -0.00041810746, -0.00026687945, -2.7334515e-06, 3.4326067e-06, -0.00028437664, -0.00026752386, -6.688769e-06, 3.2131943e-06, -0.00015109948, -0.0002650765, -1.0514272e-05, 2.9609264e-06, -1.9801768e-05, -0.00025962334, -1.4168271e-05, 2.6790735e-06, 0.00010804198, -0.00025128332, -1.7611716e-05, 2.3712018e-06, 0.00023102465, -0.00024020665, -2.0808595e-05, 2.041126e-06, 0.0003478215, -0.00022657229, -2.3726312e-05, 1.6928611e-06, 0.000457204, -0.0002105856, -2.6336e-05, 1.3305736e-06, 0.00055805227, -0.0001924754, -2.86128e-05, 9.585298e-07, 0.0006493661, -0.00017249103, -3.053608e-05, 5.8104513e-07, 0.0007302744, -0.00015089898, -3.2089603e-05, 2.0243363e-07, 0.00080004294, -0.0001279797, -3.3261647e-05, -1.7304232e-07, 0.00085808046, -0.00010402399, -3.4045068e-05, -5.412203e-07, 0.000903943, -7.932951e-05, -3.4437293e-05, -8.9808447e-07, 0.0009373362, -5.4197226e-05, -3.4440294e-05, -1.2398096e-06, 0.00095811655, -2.8927887e-05, -3.4060486e-05, -1.5628023e-06, 0.00096629, -3.8185226e-06, -3.3308566e-05, -1.8637385e-06, 0.0009620094, 2.0840904e-05, -3.219934e-05, -2.139598e-06, 0.0009455702, 4.477073e-05, -3.075146e-05, -2.3876942e-06, 0.0009174042, 6.770467e-05, -2.8987177e-05, -2.6056998e-06, 0.00087807275, 8.939263e-05, -2.6931988e-05, -2.7916674e-06, 0.00082825747, 0.00010960339, -2.461432e-05, -2.9440466e-06, 0.0007687504, 0.00012812686, -2.2065136e-05, -3.0616948e-06, 0.0007004428, 0.00014477625, -1.9317536e-05, -3.1438838e-06, 0.0006243134, 0.00015938978, -1.6406348e-05, -3.1903023e-06, 0.000541415, 0.00017183211, -1.33676895e-05, -3.2010514e-06, 0.0004528613, 0.00018199554, -1.0238536e-05, -3.1766376e-06, 0.00035981278, 0.00018980069, -7.0562724e-06, -3.1179597e-06, 0.00026346243, 0.00019519699, -3.8582616e-06, -3.0262931e-06, 0.00016502131, 0.00019816274, -6.8140974e-07, -2.9032674e-06, 6.570411e-05, 0.00019870495, 2.4382505e-06, -2.7508431e-06, -3.3284992e-05, 0.00019685866, 5.465961e-06, -2.5712827e-06, -0.0001307662, 0.00019268612, 8.368619e-06, -2.3671205e-06, -0.00022559743, 0.0001862756, 1.111513e-05, -2.1411277e-06, -0.0003166869, 0.00017773996, 1.3676734e-05, -1.896278e-06, -0.00040300505, 0.00016721482, 1.6027298e-05, -1.635709e-06, -0.00048359542, 0.00015485672, 1.814357e-05, -1.3626835e-06, -0.0005575847, 0.00014084089, 2.0005407e-05, -1.0805502e-06, -0.00062419113, 0.00012535887, 2.1595948e-05, -7.927032e-07, -0.0006827326, 0.000108616085, 2.2901751e-05, -5.025426e-07, -0.0007326324, 9.082921e-05, 2.3912902e-05, -2.1343516e-07, -0.0007734245, 7.222342e-05, 2.4623056e-05, 7.132415e-08, -0.00080475706, 5.3029675e-05, 2.502946e-05, 3.4854867e-07, -0.0008263945, 3.3481938e-05, 2.513292e-05, 6.1519495e-07, -0.0008382184, 1.3814398e-05, 2.4937726e-05, 8.6839543e-07, -0.00084022695, -5.7412394e-06, 2.445156e-05, 1.1054885e-06, -0.000832533, -2.4958403e-05, 2.3685325e-05, 1.3240457e-06, -0.0008153609, -4.36182e-05, 2.2652985e-05, 1.5218957e-06, -0.00078904204, -6.151183e-05, 2.1371345e-05, 1.6971446e-06, -0.0007540092, -7.844284e-05, 1.98598e-05, 1.8481938e-06, -0.0007107897, -9.4229166e-05, 1.8140086e-05, 1.973753e-06, -0.0006599982, -0.00010870506, 1.6235963e-05, 2.072849e-06, -0.0006023276, -0.00012172271, 1.4172929e-05, 2.1448332e-06, -0.0005385399, -0.00013315363, 1.197788e-05, 2.189382e-06, -0.0004694564, -0.0001428899, 9.678783e-06, 2.2064958e-06, -0.00039594696, -0.000150845, 7.3043298e-06, 2.1964927e-06, -0.0003189192, -0.00015695447, 4.8835964e-06, 2.16e-06, -0.00023930735, -0.00016117636, 2.4456945e-06, 2.0979417e-06, -0.000158061, -0.00016349126, 1.9438557e-08, 2.0115217e-06, -7.613381e-05, -0.00016390221, -2.3669863e-06, 1.9022065e-06, 5.5276073e-06, -0.00016243423, -4.6863383e-06, 1.7717024e-06, 8.599451e-05, -0.00015913373, -6.91262e-06, 1.6219325e-06, 0.00016436652, -0.00015406757, -9.021357e-06, 1.4550101e-06, 0.0002397816, -0.000147322, -1.09898565e-05, 1.2732113e-06, 0.00031142536, -0.00013900126, -1.2797443e-05, 1.0789458e-06, 0.00037853981, -0.00012922616, -1.4425657e-05, 8.7472654e-07, 0.0004404311, -0.000118132346, -1.585844e-05, 6.631388e-07, 0.0004964765, -0.000105868516, -1.7082273e-05, 4.4680903e-07, 0.0005461306, -9.259446e-05, -1.8086295e-05, 2.2837375e-07, 0.0005889301, -7.847905e-05, -1.8862385e-05, 1.0448686e-08, 0.00062449806, -6.369811e-05, -1.94052e-05, -2.0440125e-07, 0.00065254676, -4.84323e-05, -1.9712208e-05, -4.1369077e-07, 0.0006728795, -3.2864893e-05, -1.9783653e-05, -6.150418e-07, 0.0006853914, -1.7179666e-05, -1.9622514e-05, -8.062092e-07, 0.00069006934, -1.5587267e-06, -1.9234425e-05, -9.851045e-07, 0.00068699016, 1.3819545e-05, -1.8627563e-05, -1.1498179e-06, 0.0006763186, 2.8782508e-05, -1.7812508e-05, -1.2986367e-06, 0.00065830396, 4.316516e-05, -1.6802087e-05, -1.4300626e-06, 0.0006332757, 5.6811925e-05, -1.5611182e-05, -1.5428252e-06, 0.0006016385, 6.957828e-05, -1.4256523e-05, -1.6358925e-06, 0.000563866, 8.1332255e-05, -1.2756469e-05, -1.7084797e-06, 0.00052049453, 9.195575e-05, -1.1130761e-05, -1.7600535e-06, 0.00047211576, 0.00010134568, -9.4002735e-06, -1.7903343e-06, 0.00041936894, 0.00010941489, -7.5867533e-06, -1.7992952e-06, 0.00036293277, 0.000116092924, -5.712553e-06, -1.7871583e-06, 0.00030351683, 0.00012132655, -3.8003616e-06, -1.7543875e-06, 0.00024185305, 0.00012508009, -1.8729359e-06, -1.7016795e-06, 0.00017868665, 0.00012733552, 4.716473e-08, -1.6299514e-06, 0.00011476754, 0.00012809242, 1.9378356e-06, -1.540327e-06, 5.0841467e-05, 0.0001273677, 3.7776758e-06, -1.43412e-06, -1.2358492e-05, 0.00012519505, 5.5462247e-06, -1.3128151e-06, -7.412017e-05, 0.000121624274, 7.224183e-06, -1.1780489e-06, -0.0001337602, 0.00011672055, 8.793616e-06, -1.0315878e-06, -0.00019063136, 0.00011056328, 1.0238141e-05, -8.753053e-07, -0.00024412952, 0.00010324503, 1.154309e-05, -7.1115886e-07, -0.00029369982, 9.487021e-05, 1.269565e-05, -5.4116543e-07, -0.00033884228, 8.555365e-05, 1.3684982e-05, -3.673775e-07, -0.00037911665, 7.541913e-05, 1.4502314e-05, -1.918583e-07, -0.00041414646, 6.459776e-05, 1.5141006e-05, -1.6657985e-08, -0.00044362227, 5.322641e-05, 1.5596595e-05, 1.5621004e-07, -0.00046730423, 4.1445935e-05, 1.5866808e-05, 3.2479178e-07, -0.00048502345, 2.9399558e-05, 1.5951551e-05, 4.872143e-07, -0.000496683, 1.7231143e-05, 1.5852878e-05, 6.417063e-07, -0.00050225767, 5.0835165e-06, 1.5574926e-05, 7.866165e-07, -0.000501793, -6.9031535e-06, 1.5123837e-05, 9.204313e-07, -0.00049540366, -1.8592944e-05, 1.4507653e-05, 1.0417896e-06, -0.00048327097, -2.985567e-05, 1.37361885e-05, 1.1494964e-06, -0.00046563946, -4.0568302e-05, 1.2820891e-05, 1.2425335e-06, -0.00044281324, -5.061626e-05, 1.17746795e-05, 1.3200689e-06, -0.00041515133, -5.989461e-05, 1.0611769e-05, 1.3814628e-06, -0.00038306252, -6.830909e-05, 9.347489e-06, 1.4262722e-06, -0.00034699994, -7.5777054e-05, 7.998085e-06, 1.4542526e-06, -0.00030745493, -8.22282e-05, 6.580511e-06, 1.4653576e-06, -0.0002649508, -8.760522e-05, 5.1122324e-06, 1.4597363e-06, -0.00022003613, -9.186418e-05, 3.6110046e-06, 1.437728e-06, -0.00017327811, -9.4974865e-05, 2.0946684e-06, 1.3998554e-06, -0.00012525555, -9.692086e-05, 5.8094145e-07, 1.3468156e-06, -7.655202e-05, -9.769953e-05, -9.127852e-07, 1.2794687e-06, -2.7749007e-05, -9.732179e-05, -2.3696427e-06, 1.198826e-06, 2.058078e-05, -9.581178e-05, -3.7734703e-06, 1.1060347e-06, 6.7879904e-05, -9.320637e-05, -5.1089905e-06, 1.0023633e-06, 0.000113612405, -8.955446e-05, -6.3619723e-06, 8.8918443e-07, 0.00015726963, -8.491628e-05, -7.5193757e-06, 7.6795754e-07, 0.00019837571, -7.9362464e-05, -8.569485e-06, 6.402103e-07, 0.00023649246, -7.2973075e-05, -9.502019e-06, 5.075201e-07, 0.00027122386, -6.5836495e-05, -1.0308231e-05, 3.7149482e-07, 0.00030221997, -5.8048292e-05, -1.0980981e-05, 2.3375374e-07, 0.0003291801, -4.970997e-05, -1.1514789e-05, 9.590874e-08, 0.0003518556, -4.09277e-05, -1.1905875e-05, -4.045425e-08, 0.0003700517, -3.1811025e-05, -1.2152172e-05, -1.7379317e-07, 0.0003836291, -2.247151e-05, -1.2253321e-05, -3.026269e-07, 0.00039250444, -1.3021434e-05, -1.2210649e-05, -4.2555126e-07, 0.00039665043, -3.5724718e-06, -1.2027122e-05, -5.4125417e-07, 0.00039609513, 5.7655866e-06, -1.1707282e-05, -6.48529e-07, 0.00039092085, 1.488608e-05, -1.1257177e-05, -7.46287e-07, 0.00038126216, 2.3686656e-05, -1.06842535e-05, -8.3356764e-07, 0.00036730347, 3.2070388e-05, -9.997255e-06, -9.095478e-07, 0.00034927618, 3.99468e-05, -9.206096e-06, -9.735488e-07, 0.00032745497, 4.7232814e-05, -8.32173e-06, -1.0250419e-06, 0.00030215413, 5.3853582e-05, -7.3560022e-06, -1.0636519e-06, 0.00027372318, 5.9743223e-05, -6.3214984e-06, -1.0891589e-06, 0.00024254216, 6.484542e-05, -5.231389e-06, -1.1014981e-06, 0.00020901674, 6.911395e-05, -4.0992645e-06, -1.1007583e-06, 0.00017357318, 7.2512994e-05, -2.9389716e-06, -1.0871773e-06, 0.00013665296, 7.501741e-05, -1.7644494e-06, -1.0611384e-06, 9.87074e-05, 7.6612865e-05, -5.895656e-07, -1.0231615e-06, 6.0192346e-05, 7.729579e-05, 5.720419e-07, -9.738964e-07, 2.1562724e-05, 7.707322e-05, 1.70712e-06, -9.141121e-07, -1.6732654e-05, 7.596262e-05, 2.802946e-06, -8.446863e-07, -5.425622e-05, 7.399141e-05, 3.8474677e-06, -7.6659353e-07, -9.058652e-05, 7.119654e-05, 4.82943e-06, -6.808917e-07, -0.00012532285, 6.762388e-05, 5.7384927e-06, -5.887091e-07, -0.0001580895, 6.332756e-05, 6.565335e-06, -4.912297e-07, -0.00018853977, 5.8369184e-05, 7.3017445e-06, -3.8967877e-07, -0.00021635942, 5.2817e-05, 7.940697e-06, -2.8530778e-07, -0.00024126982, 4.6744997e-05, 8.476415e-06, -1.7937968e-07, -0.00026303058, 4.0231964e-05, 8.904414e-06, -7.3153934e-08, -0.00028144172, 3.3360477e-05, 9.221534e-06, 3.2127932e-08, -0.00029634527, 2.6215896e-05, 9.425953e-06, 1.3525641e-07, -0.00030762635, 1.8885325e-05, 9.517186e-06, 2.350675e-07, -0.00031521395, 1.1456575e-05, 9.496067e-06, 3.3045538e-07, -0.0003190809, 4.017131e-06, 9.3647195e-06, 4.2038428e-07, -0.00031924344, -3.3468475e-06, 9.126507e-06, 5.038993e-07, -0.00031576038, -1.0551507e-05, 8.785978e-06, 5.80136e-07, -0.00030873172, -1.7516233e-05, 8.348788e-06, 6.48329e-07, -0.00029829674, -2.4164523e-05, 7.821619e-06, 7.0781925e-07, -0.00028463174, -3.042481e-05, 7.2120833e-06, 7.580597e-07, -0.00026794747, -3.6231206e-05, 6.5286226e-06, 7.9861974e-07, -0.00024848603, -4.152417e-05, 5.7803913e-06, 8.291885e-07, -0.0002265176, -4.625109e-05, 4.9771434e-06, 8.4957605e-07, -0.0002023368, -5.036678e-05, 4.1291064e-06, 8.597141e-07, -0.00017625892, -5.383387e-05, 3.2468565e-06, 8.59654e-07, -0.00014861595, -5.6623125e-05, 2.3411897e-06, 8.4956497e-07, -0.00011975233, -5.8713624e-05, 1.4229928e-06, 8.2972946e-07, -9.002095e-05, -6.0092883e-05, 5.031167e-07, 8.005384e-07, -5.977878e-05, -6.0756858e-05, -4.0774938e-07, 7.624847e-07, -2.9382736e-05, -6.0709834e-05, -1.2991989e-06, 7.161559e-07, 8.14462e-07, -5.9964248e-05, -2.1612236e-06, 6.622257e-07, 3.0468289e-05, -5.8540416e-05, -2.9843227e-06, 6.0144475e-07, 5.9246275e-05, -5.6466146e-05, -3.7596046e-06, 5.346306e-07, 8.6831635e-05, -5.377632e-05, -4.4788794e-06, 4.6265728e-07, 0.000112926675, -5.0512335e-05, -5.1347433e-06, 3.86444e-07, 0.00013725593, -4.6721547e-05, -5.7206485e-06, 3.0694392e-07, 0.00015956897, -4.2456617e-05, -6.230967e-06, 2.2513252e-07, 0.00017964284, -3.777479e-05, -6.6610396e-06, 1.4199584e-07, 0.00019728423, -3.2737193e-05, -7.0072147e-06, 5.8518935e-08, 0.0002123312, -2.7408027e-05, -7.2668718e-06, -2.4325521e-08, 0.00022465452, -2.1853803e-05, -7.438435e-06, -1.0558829e-07, 0.00023415861, -1.6142507e-05, -7.5213766e-06, -1.8435419e-07, 0.00024078209, -1.0342813e-05, -7.516201e-06, -2.597521e-07, 0.0002444979, -4.523257e-06, -7.4244263e-06, -3.3096438e-07, 0.0002453131, 1.2485418e-06, -7.2485464e-06, -3.9723534e-07, 0.00024326815, 6.9066514e-06, -6.991987e-06, -4.5787905e-07, 0.00023843585, 1.2387563e-05, -6.6590515e-06, -5.1228614e-07, 0.00023092006, 1.7630884e-05, -6.2548543e-06, -5.599294e-07, 0.0002208539, 2.2579985e-05, -5.7852503e-06, -6.0036876e-07, 0.00020839775, 2.718259e-05, -5.256753e-06, -6.3325484e-07, 0.0001937369, 3.139131e-05, -4.676449e-06, -6.583313e-07, 0.00017707904, 3.516412e-05, -4.051906e-06, -6.754366e-07, 0.00015865147, 3.846473e-05, -3.3910783e-06, -6.84504e-07, 0.00013869806, 4.1262923e-05, -2.702206e-06, -6.8556096e-07, 0.00011747629, 4.3534823e-05, -1.9937172e-06, -6.78727e-07, 9.5253905e-05, 4.526303e-05, -1.274126e-06, -6.642111e-07, 7.2305746e-05, 4.6436733e-05, -5.5193306e-07, -6.423075e-07, 4.891038e-05, 4.705172e-05, 1.6447315e-07, -6.133911e-07, 2.5346864e-05, 4.7110312e-05, 8.6691074e-07, -5.779116e-07, 1.8914722e-06, 4.662124e-05, 1.5474963e-06, -5.363872e-07, -2.1185442e-05, 4.559942e-05, 2.1987307e-06, -4.893973e-07, -4.3622476e-05, 4.4065688e-05, 2.81358e-06, -4.375749e-07, -6.517005e-05, 4.204645e-05, 3.3855483e-06, -3.815984e-07, -8.55931e-05, 3.9573297e-05, 3.9087445e-06, -3.2218284e-07, -0.00010467357, 3.668254e-05, 4.37794e-06, -2.6007118e-07, -0.00012221262, 3.341471e-05, 4.788619e-06, -1.9602507e-07, -0.00013803263, 2.9814035e-05, 5.137018e-06, -1.3081595e-07, -0.00015197888, 2.5927835e-05, 5.420156e-06, -6.521575e-08, -0.000163921, 2.1805956e-05, 5.6358576e-06, 1.1952672e-11, -0.000173754, 1.7500131e-05, 5.7827638e-06, 6.4120634e-08, -0.00018139913, 1.3063353e-05, 5.860334e-06, 1.263892e-07, -0.0001868043, 8.549245e-06, 5.8688393e-06, 1.8612985e-07, -0.00018994427, 4.011421e-06, 5.8093447e-06, 2.4269556e-07, -0.00019082046, -4.971275e-07, 5.683684e-06, 2.9548684e-07, -0.00018946052, -4.924638e-06, 5.494426e-06, 3.4395785e-07, -0.00018591754, -9.221154e-06, 5.2448327e-06, 3.8762184e-07, -0.00018026902, -1.3339076e-05, 4.9388077e-06, 4.2605583e-07, -0.0001726156, -1.7233668e-05, 4.580844e-06, 4.589044e-07, -0.00016307941, -2.0863534e-05, 4.1759586e-06, 4.8588265e-07, -0.00015180242, -2.4191033e-05, 3.7296281e-06, 5.0677835e-07, -0.00013894434, -2.7182663e-05, 3.2477167e-06, 5.214532e-07, -0.00012468056, -2.9809366e-05, 2.7364015e-06, 5.2984313e-07, -0.00010919985, -3.2046803e-05, 2.202096e-06, 5.319579e-07, -9.27019e-05, -3.3875545e-05, 1.651373e-06, 5.278795e-07, -7.5394855e-05, -3.5281228e-05, 1.090884e-06, 5.177603e-07, -5.7492776e-05, -3.625462e-05, 5.272819e-07, 5.018201e-07, -3.921303e-05, -3.679166e-05, -3.285569e-08, 4.803421e-07, -2.0773752e-05, -3.6893394e-05, -5.83102e-07, 4.5366892e-07, -2.3912733e-06, -3.6565907e-05, -1.1172526e-06, 4.221975e-07, 1.5722333e-05, -3.5820143e-05, -1.6293935e-06, 3.8637359e-07, 3.336164e-05, -3.4671713e-05, -2.113965e-06, 3.466858e-07, 5.033014e-05, -3.3140623e-05, -2.5658196e-06, 3.0365925e-07, 6.644237e-05, -3.1250976e-05, -2.9802754e-06, 2.5784885e-07, 8.152586e-05, -2.9030636e-05, -3.3531614e-06, 2.0983232e-07, 9.542295e-05, -2.6510814e-05, -3.6808583e-06, 1.6020327e-07, 0.00010799231, -2.3725677e-05, -3.960331e-06, 1.0956389e-07, 0.00011911037, -2.0711894e-05, -4.189153e-06, 5.8517998e-08, 0.0001286724, -1.750816e-05, -4.365525e-06, 7.663899e-09, 0.00013659344, -1.41547325e-05, -4.488286e-06, -4.2412374e-08, 0.00014280893, -1.0692924e-05, -4.556914e-06, -9.114367e-08, 0.00014727515, -7.1646145e-06, -4.5715233e-06, -1.3798794e-07, 0.00014996933, -3.6117533e-06, -4.5328516e-06, -1.8243412e-07, 0.00015088962, -7.587294e-08, -4.4422413e-06, -2.2400754e-07, 0.00015005471, 3.4023838e-06, -4.301613e-06, -2.622747e-07, 0.0001475033, 6.7837195e-06, -4.1134344e-06, -2.968478e-07, 0.00014329332, 1.0030616e-05, -3.880684e-06, -3.2738822e-07, 0.00013750092, 1.3107738e-05, -3.6068036e-06, -3.536098e-07, 0.00013021928, 1.5982303e-05, -3.2956561e-06, -3.752812e-07, 0.00012155731, 1.8624423e-05, -2.9514704e-06, -3.9222766e-07, 0.00011163802, 2.1007401e-05, -2.5787865e-06, -4.043321e-07, 0.00010059696, 2.3107985e-05, -2.182399e-06, -4.1153544e-07, 8.8580375e-05, 2.4906572e-05, -1.7672962e-06, -4.138364e-07, 7.574336e-05, 2.6387395e-05, -1.3386002e-06, -4.1129053e-07, 6.2247935e-05, 2.7538621e-05, -9.0150434e-07, -4.0400852e-07, 4.826102e-05, 2.8352426e-05, -4.6121215e-07, -3.9215408e-07, 3.395243e-05, 2.8825028e-05, -2.2877371e-08, -3.759412e-07, 1.9492882e-05, 2.8956656e-05, 4.0845538e-07, -3.5563068e-07, 5.0519816e-06, 2.8751478e-05, 8.279069e-07, -3.315265e-07, -9.203712e-06, 2.8217493e-05, 1.2308172e-06, -3.0397143e-07, -2.3112565e-05, 2.7366372e-05, 1.6127958e-06, -2.7334247e-07, -3.6519654e-05, 2.6213258e-05, 1.9697682e-06, -2.4004595e-07, -4.9278453e-05, 2.4776538e-05, 2.298017e-06, -2.045123e-07, -6.125238e-05, 2.3077575e-05, 2.5942204e-06, -1.6719062e-07, -7.2316216e-05, 2.1140404e-05, 2.8554823e-06, -1.2854323e-07, -8.2357365e-05, 1.8991419e-05, 3.0793606e-06, -8.904007e-08, -9.127695e-05, 1.6659023e-05, 3.2638857e-06, -4.9153147e-08, -9.899071e-05, 1.4173269e-05, 3.4075777e-06, -9.350997e-09, -0.00010542977, 1.1565476e-05, 3.509453e-06, 2.9906634e-08, -0.000110541114, 8.8678535e-06, 3.5690296e-06, 6.8173996e-08, -0.000114288, 6.113115e-06, 3.5863227e-06, 1.05024256e-07, -0.00011665008, 3.3340827e-06, 3.561837e-06, 1.4005413e-07, -0.00011762337, 5.6331345e-07, 3.4965524e-06, 1.7288812e-07, -0.000117220006, -2.1672777e-06, 3.3919043e-06, 2.0318245e-07};
endpackage
`endif
