`ifndef COEFFICIENTS_FX_SV_
`define COEFFICIENTS_FX_SV_
package Coefficients_Fx;
	localparam N = 4;
	localparam M = 4;
	localparam COEFF_BIAS = 48;
	localparam logic signed[63:0] Lfr[0:3] = {64'd279614656416265, 64'd279614656416265, 64'd277224080786690, 64'd277224080786690};
	localparam logic signed[63:0] Lfi[0:3] = {64'd8476895612029, - 64'd8476895612029, 64'd3418304876175, - 64'd3418304876175};
	localparam logic signed[63:0] Lbr[0:3] = {64'd279614656416265, 64'd279614656416265, 64'd277224080786690, 64'd277224080786690};
	localparam logic signed[63:0] Lbi[0:3] = {64'd8476895612029, - 64'd8476895612029, 64'd3418304876175, - 64'd3418304876175};
	localparam logic signed[63:0] Wfr[0:3] = {64'd568700833, 64'd568700833, 64'd169265178, 64'd169265178};
	localparam logic signed[63:0] Wfi[0:3] = {64'd21481769, - 64'd21481769, 64'd325649128, - 64'd325649128};
	localparam logic signed[63:0] Wbr[0:3] = {- 64'd568700833, - 64'd568700833, - 64'd169265178, - 64'd169265178};
	localparam logic signed[63:0] Wbi[0:3] = {- 64'd21481769, 64'd21481769, - 64'd325649128, 64'd325649128};
	localparam logic signed[63:0] Ffr[0:3][0:99] = '{
		'{64'd209367917907850816, 64'd12940596353402938, - 64'd896381733843701, 64'd5773941780322, 64'd215697698286196160, 64'd12377665357757680, - 64'd899926540939321, 64'd6975477820499, 64'd221744772881992928, 64'd11809873366082668, - 64'd902572342792447, 64'd8155642492392, 64'd227506861175543360, 64'd11237819785294670, - 64'd904327652903445, 64'd9313576045912, 64'd232981981547220352, 64'd10662100720251796, - 64'd905201726880791, 64'd10448450412235, 64'd238168449494480192, 64'd10083308447572872, - 64'd905204544538224, 64'd11559469602358, 64'd243064875588293056, 64'd9502030899551228, - 64'd904346791523053, 64'd12645870070256, 64'd247670163174130496, 64'd8918851158529572, - 64'd902639840498836, 64'd13706921040752, 64'd251983505822829600, 64'd8334346962088413, - 64'd900095731905798, 64'd14741924802207, 64'd256004384536825024, 64'd7749090219385679, - 64'd896727154322443, 64'd15750216964190, 64'd259732564717406848, 64'd7163646538970562, - 64'd892547424451934, 64'd16731166680303, 64'd263168092898817728, 64'd6578574768379709, - 64'd887570466756864, 64'd17684176836396, 64'd266311293255155840, 64'd5994426545808893, - 64'd881810792766088, 64'd18608684204390, 64'd269162763886189760, 64'd5411745864138234, - 64'd875283480077328, 64'd19504159562015, 64'd271723372888330976, 64'd4831068647573912, - 64'd868004151079220, 64'd20370107778738, 64'd273994254217131520, 64'd4252922341153986, - 64'd859988951416491, 64'd21206067868235, 64'd275976803347800640, 64'd3677825513350828, - 64'd851254528221888, 64'd22011613007759, 64'd277672672740341760, 64'd3106287471987255, - 64'd841818008138399, 64'd22786350524788, 64'd279083767116018560, 64'd2538807893668153, - 64'd831696975155255, 64'd23529921851380, 64'd280212238551954656, 64'd1975876466914083, - 64'd820909448281046, 64'd24242002446658, 64'd281060481400761920, 64'd1417972549168047, - 64'd809473859077193, 64'd24922301687903, 64'd281631127042172608, 64'd865564837831255, - 64'd797409029074828, 64'd25570562730737, 64'd281927038473727296, 64'd319111055468575, - 64'd784734147098001, 64'd26186562338910, 64'd281951304747633280, - 64'd220942350690998, - 64'd771468746515904, 64'd26770110684226, 64'd281707235260971136, - 64'd754160494848410, - 64'd757632682446620, 64'd27321051117161},
		'{64'd209367917907958112, 64'd12940596353398758, - 64'd896381733843569, 64'd5773941780326, 64'd215697698286299968, 64'd12377665357753640, - 64'd899926540939193, 64'd6975477820503, 64'd221744772882093280, 64'd11809873366078768, - 64'd902572342792324, 64'd8155642492396, 64'd227506861175640128, 64'd11237819785290916, - 64'd904327652903325, 64'd9313576045915, 64'd232981981547313472, 64'd10662100720248186, - 64'd905201726880675, 64'd10448450412239, 64'd238168449494569664, 64'd10083308447569412, - 64'd905204544538113, 64'd11559469602361, 64'd243064875588378848, 64'd9502030899547916, - 64'd904346791522946, 64'd12645870070259, 64'd247670163174212544, 64'd8918851158526408, - 64'd902639840498734, 64'd13706921040755, 64'd251983505822907872, 64'd8334346962085402, - 64'd900095731905700, 64'd14741924802210, 64'd256004384536899488, 64'd7749090219382820, - 64'd896727154322349, 64'd15750216964192, 64'd259732564717477504, 64'd7163646538967858, - 64'd892547424451845, 64'd16731166680306, 64'd263168092898884544, 64'd6578574768377158, - 64'd887570466756779, 64'd17684176836398, 64'd266311293255218816, 64'd5994426545806495, - 64'd881810792766008, 64'd18608684204392, 64'd269162763886248896, 64'd5411745864135991, - 64'd875283480077252, 64'd19504159562017, 64'd271723372888386208, 64'd4831068647571824, - 64'd868004151079148, 64'd20370107778739, 64'd273994254217182848, 64'd4252922341152053, - 64'd859988951416425, 64'd21206067868237, 64'd275976803347848064, 64'd3677825513349051, - 64'd851254528221826, 64'd22011613007760, 64'd277672672740385280, 64'd3106287471985634, - 64'd841818008138342, 64'd22786350524789, 64'd279083767116058240, 64'd2538807893666684, - 64'd831696975155202, 64'd23529921851382, 64'd280212238551990528, 64'd1975876466912769, - 64'd820909448280998, 64'd24242002446659, 64'd281060481400793856, 64'd1417972549166887, - 64'd809473859077149, 64'd24922301687904, 64'd281631127042200768, 64'd865564837830247, - 64'd797409029074788, 64'd25570562730738, 64'd281927038473751616, 64'd319111055467717, - 64'd784734147097966, 64'd26186562338911, 64'd281951304747653824, - 64'd220942350691705, - 64'd771468746515874, 64'd26770110684226, 64'd281707235260987936, - 64'd754160494848966, - 64'd757632682446594, 64'd27321051117161},
		'{64'd208807812964745760, 64'd12908849052433810, - 64'd876670745151696, 64'd74765294786063, 64'd215125675568580832, 64'd12364546145487408, - 64'd846574522093956, 64'd73015021252188, 64'd221174290868974432, 64'd11831835552141554, - 64'd817058095947687, 64'd71289534886562, 64'd226959418591712288, 64'd11310571551516128, - 64'd788115257212276, 64'd69588744339475, 64'd232486745611835648, 64'd10800608470538784, - 64'd759739766193057, 64'd67912551711317, 64'd237761885990934528, 64'd10301800737227882, - 64'd731925356245339, 64'd66260852784717, 64'd242790381040674016, 64'd9814002932348062, - 64'd704665736931800, 64'd64633537252140, 64'd247577699411748000, 64'd9337069839467642, - 64'd677954597094628, 64'd63030488938973, 64'd252129237207467552, 64'd8870856493446672, - 64'd651785607843809, 64'd61451586022165, 64'd256450318121207584, 64'd8415218227384312, - 64'd626152425462938, 64'd59896701244465, 64'd260546193596947328, 64'd7970010718053768, - 64'd601048694233914, 64'd58365702124314, 64'd264422043012156608, 64'd7535090029852914, - 64'd576468049181897, 64'd56858451161428, 64'd268082973882291328, 64'd7110312657298326, - 64'd552404118741850, 64'd55374806038149, 64'd271534022086178720, 64'd6695535566090250, - 64'd528850527348025, 64'd53914619816584, 64'd274780152111582368, 64'd6290616232775662, - 64'd505800897947707, 64'd52477741131608, 64'd277826257320254464, 64'd5895412683036402, - 64'd483248854440530, 64'd51064014379769, 64'd280677160231793856, 64'd5509783528628952, - 64'd461188024044683, 64'd49673279904155, 64'd283337612825642464, 64'd5133588003002269, - 64'd439612039591281, 64'd48305374175258, 64'd285812296860565440, 64'd4766685995619665, - 64'd418514541748187, 64'd46960129967909, 64'd288105824210973600, 64'd4408938085010547, - 64'd397889181174568, 64'd45637376534320, 64'd290222737219459648, 64'd4060205570577469, - 64'd377729620607419, 64'd44336939773278, 64'd292167509064932096, 64'd3720350503183700, - 64'd358029536881318, 64'd43058642395570, 64'd293944544145742976, 64'd3389235714546153, - 64'd338782622882642, 64'd41802304085651, 64'd295558178477218880, 64'd3066724845458330, - 64'd319982589439454, 64'd40567741659640, 64'd297012680103015168, 64'd2752682372867516, - 64'd301623167148285, 64'd39354769219676},
		'{64'd208807812965074720, 64'd12908849052420436, - 64'd876670745151279, 64'd74765294786075, 64'd215125675568903712, 64'd12364546145474280, - 64'd846574522093546, 64'd73015021252200, 64'd221174290869291296, 64'd11831835552128672, - 64'd817058095947284, 64'd71289534886574, 64'd226959418592023200, 64'd11310571551503488, - 64'd788115257211881, 64'd69588744339487, 64'd232486745612140672, 64'd10800608470526384, - 64'd759739766192669, 64'd67912551711329, 64'd237761885991233696, 64'd10301800737215720, - 64'd731925356244959, 64'd66260852784729, 64'd242790381040967424, 64'd9814002932336134, - 64'd704665736931427, 64'd64633537252152, 64'd247577699412035712, 64'd9337069839455944, - 64'd677954597094262, 64'd63030488938984, 64'd252129237207749632, 64'd8870856493435206, - 64'd651785607843450, 64'd61451586022176, 64'd256450318121484064, 64'd8415218227373072, - 64'd626152425462585, 64'd59896701244476, 64'd260546193597218304, 64'd7970010718042754, - 64'd601048694233569, 64'd58365702124324, 64'd264422043012422080, 64'd7535090029842121, - 64'd576468049181558, 64'd56858451161439, 64'd268082973882551424, 64'd7110312657287754, - 64'd552404118741518, 64'd55374806038159, 64'd271534022086433504, 64'd6695535566079894, - 64'd528850527347700, 64'd53914619816594, 64'd274780152111831872, 64'd6290616232765520, - 64'd505800897947388, 64'd52477741131617, 64'd277826257320498752, 64'd5895412683026470, - 64'd483248854440218, 64'd51064014379779, 64'd280677160232033024, 64'd5509783528619232, - 64'd461188024044378, 64'd49673279904164, 64'd283337612825876544, 64'd5133588002992756, - 64'd439612039590981, 64'd48305374175267, 64'd285812296860794496, 64'd4766685995610355, - 64'd418514541747894, 64'd46960129967918, 64'd288105824211197728, 64'd4408938085001438, - 64'd397889181174281, 64'd45637376534328, 64'd290222737219678848, 64'd4060205570568558, - 64'd377729620607138, 64'd44336939773286, 64'd292167509065146496, 64'd3720350503174987, - 64'd358029536881044, 64'd43058642395578, 64'd293944544145952640, 64'd3389235714537633, - 64'd338782622882373, 64'd41802304085659, 64'd295558178477423808, 64'd3066724845450001, - 64'd319982589439191, 64'd40567741659648, 64'd297012680103215488, 64'd2752682372859375, - 64'd301623167148028, 64'd39354769219683}};
	localparam logic signed[63:0] Ffi[0:3][0:99] = '{
		'{- 64'd256127510662709344, 64'd15852187053065382, 64'd314423079823242, - 64'd41164091899801, - 64'd248129395814423328, 64'd16137135790239808, 64'd285349582355099, - 64'd40718142853921, - 64'd239993514431440960, 64'd16403248028101054, 64'd256361481670483, - 64'd40238955728992, - 64'd231729291000865696, 64'd16650501866890788, 64'd227485287792818, - 64'd39727393821403, - 64'd223346156401711360, 64'd16878893603318750, 64'd198747079143438, - 64'd39184340614075, - 64'd214853538860987136, 64'd17088437510854180, 64'd170172483044807, - 64'd38610698688936, - 64'd206260855023252512, 64'd17279165605622898, 64'd141786656891765, - 64'd38007388634573, - 64'd197577501140738400, 64'd17451127398309160, 64'd113614270000494, - 64'd37375347950170, - 64'd188812844390932416, 64'd17604389632469850, 64'd85679486144150, - 64'd36715529946819, - 64'd179976214328316672, 64'd17739036009676462, 64'd58005946783340, - 64'd36028902647275, - 64'd171076894476740416, 64'd17855166901907766, 64'd30616754998861, - 64'd35316447685221, - 64'd162124114068693760, 64'd17952899051622972, 64'd3534460133363, - 64'd34579159205100, - 64'd153127039937533984, 64'd18032365259951640, - 64'd23218956852172, - 64'd33818042763551, - 64'd144094768568495984, 64'd18093714063442580, - 64'd49622097301960, - 64'd33034114233470, - 64'd135036318314095360, 64'd18137109399819340, - 64'd75654158064577, - 64'd32228398711708, - 64'd125960621779307344, 64'd18162730263194952, - 64'd101294943964075, - 64'd31401929431406, - 64'd116876518381679152, 64'd18170770349202968, - 64'd126524879540126, - 64'd30555746679929, - 64'd107792747091301296, 64'd18161437690505888, - 64'd151325020055019, - 64'd29690896723379, - 64'd98717939355333744, 64'd18134954283145528, - 64'd175677061766010, - 64'd28808430738610, - 64'd89660612211549136, 64'd18091555704202836, - 64'd199563351462307, - 64'd27909403753678, - 64'd80629161595120784, 64'd18031490721237340, - 64'd222966895266617, - 64'd26994873597632, - 64'd71631855842647376, 64'd17955020893978248, - 64'd245871366701920, - 64'd26065899860521, - 64'd62676829397171616, 64'd17862420168741000, - 64'd268261114024824, - 64'd25123542864488, - 64'd53772076717708672, 64'd17753974466044040, - 64'd290121166827504, - 64'd24168862646791, - 64'd44925446396568800, 64'd17629981261901270, - 64'd311437241910954, - 64'd23202917955564},
		'{64'd256127510662618048, - 64'd15852187053061658, - 64'd314423079823345, 64'd41164091899796, 64'd248129395814329408, - 64'd16137135790235982, - 64'd285349582355205, 64'd40718142853917, 64'd239993514431344512, - 64'd16403248028097132, - 64'd256361481670592, 64'd40238955728987, 64'd231729291000766880, - 64'd16650501866886776, - 64'd227485287792931, 64'd39727393821398, 64'd223346156401610272, - 64'd16878893603314652, - 64'd198747079143554, 64'd39184340614070, 64'd214853538860883936, - 64'd17088437510849998, - 64'd170172483044925, 64'd38610698688932, 64'd206260855023147264, - 64'd17279165605618642, - 64'd141786656891886, 64'd38007388634568, 64'd197577501140631296, - 64'd17451127398304828, - 64'd113614270000618, 64'd37375347950165, 64'd188812844390823520, - 64'd17604389632465452, - 64'd85679486144276, 64'd36715529946814, 64'd179976214328206144, - 64'd17739036009672002, - 64'd58005946783468, 64'd36028902647270, 64'd171076894476628416, - 64'd17855166901903252, - 64'd30616754998991, 64'd35316447685216, 64'd162124114068580352, - 64'd17952899051618404, - 64'd3534460133494, 64'd34579159205095, 64'd153127039937419296, - 64'd18032365259947028, 64'd23218956852039, 64'd33818042763546, 64'd144094768568380176, - 64'd18093714063437924, 64'd49622097301825, 64'd33034114233465, 64'd135036318313978528, - 64'd18137109399814648, 64'd75654158064441, 64'd32228398711703, 64'd125960621779189600, - 64'd18162730263190228, 64'd101294943963937, 64'd31401929431400, 64'd116876518381560656, - 64'd18170770349198216, 64'd126524879539988, 64'd30555746679924, 64'd107792747091182144, - 64'd18161437690501116, 64'd151325020054879, 64'd29690896723374, 64'd98717939355214080, - 64'd18134954283140736, 64'd175677061765869, 64'd28808430738604, 64'd89660612211429088, - 64'd18091555704198032, 64'd199563351462166, 64'd27909403753672, 64'd80629161595000416, - 64'd18031490721232532, 64'd222966895266475, 64'd26994873597627, 64'd71631855842526880, - 64'd17955020893973436, 64'd245871366701779, 64'd26065899860516, 64'd62676829397051056, - 64'd17862420168736188, 64'd268261114024682, 64'd25123542864483, 64'd53772076717588176, - 64'd17753974466039234, 64'd290121166827362, 64'd24168862646785, 64'd44925446396448464, - 64'd17629981261896476, 64'd311437241910812, 64'd23202917955559},
		'{- 64'd779901327374593024, 64'd28766736086525376, - 64'd1388026451385535, 64'd51147782792348, - 64'd765587272939073280, 64'd28489063021489052, - 64'd1377710692110832, 64'd51283306989880, - 64'd751412666690274560, 64'd28208973279885160, - 64'd1367185227349448, 64'd51395528697467, - 64'd737378672460398336, 64'd27926644138938352, - 64'd1356460265322528, 64'd51485100856128, - 64'd723486366557601280, 64'd27642248428922260, - 64'd1345545784674669, 64'd51552665436647, - 64'd709736739972521728, 64'd27355954600898964, - 64'd1334451537574361, 64'd51598853525713, - 64'd696130700551027584, 64'd27067926794082408, - 64'd1323187052806982, 64'd51624285413561, - 64'd682669075133381504, 64'd26778324902811884, - 64'd1311761638859439, 64'd51629570683067, - 64'd669352611660017792, 64'd26487304643121916, - 64'd1300184386995524, 64'd51615308300201, - 64'd656181981244139648, 64'd26195017618895720, - 64'd1288464174321125, 64'd51582086705768, - 64'd643157780211344768, 64'd25901611387589656, - 64'd1276609666838425, 64'd51530483908368, - 64'd630280532106499840, 64'd25607229525516912, - 64'd1264629322488288, 64'd51461067578499, - 64'd617550689668085120, 64'd25312011692679012, - 64'd1252531394180023, 64'd51374395143739, - 64'd604968636770238464, 64'd25016093697134284, - 64'd1240323932807792, 64'd51271013884931, - 64'd592534690332733568, 64'd24719607558892892, - 64'd1228014790252892, 64'd51151461033313, - 64'd580249102199129728, 64'd24422681573328616, - 64'd1215611622371236, 64'd51016263868523, - 64'd568112060983341312, 64'd24125440374097968, - 64'd1203121891965334, 64'd50865939817420, - 64'd556123693884869504, 64'd23828004995557668, - 64'd1190552871740133, 64'd50700996553656, - 64'd544284068472954624, 64'd23530492934672044, - 64'd1177911647242071, 64'd50521932097940, - 64'd532593194439903232, 64'd23233018212402304, - 64'd1165205119780762, 64'd50329234918942, - 64'd521051025323850944, 64'd22935691434570068, - 64'd1152440009332711, 64'd50123384034762, - 64'd509657460201228672, 64'd22638619852188048, - 64'd1139622857426528, 64'd49904849114941, - 64'd498412345349195520, 64'd22341907421251000, - 64'd1126760030009089, 64'd49674090582920, - 64'd487315475878314432, 64'd22045654861980704, - 64'd1113857720292146, 64'd49431559718926, - 64'd476366597335741120, 64'd21749959717518912, - 64'd1100921951578898, 64'd49177698763224},
		'{64'd779901327374501888, - 64'd28766736086521656, 64'd1388026451385433, - 64'd51147782792353, 64'd765587272938979456, - 64'd28489063021485228, 64'd1377710692110726, - 64'd51283306989884, 64'd751412666690178304, - 64'd28208973279881232, 64'd1367185227349340, - 64'd51395528697472, 64'd737378672460299648, - 64'd27926644138934324, 64'd1356460265322416, - 64'd51485100856132, 64'd723486366557500416, - 64'd27642248428918144, 64'd1345545784674554, - 64'd51552665436652, 64'd709736739972418560, - 64'd27355954600894760, 64'd1334451537574243, - 64'd51598853525718, 64'd696130700550922368, - 64'd27067926794078116, 64'd1323187052806861, - 64'd51624285413566, 64'd682669075133274368, - 64'd26778324902807512, 64'd1311761638859315, - 64'd51629570683072, 64'd669352611659908864, - 64'd26487304643117472, 64'd1300184386995398, - 64'd51615308300206, 64'd656181981244028800, - 64'd26195017618891204, 64'd1288464174320996, - 64'd51582086705773, 64'd643157780211232128, - 64'd25901611387585068, 64'd1276609666838294, - 64'd51530483908373, 64'd630280532106385792, - 64'd25607229525512260, 64'd1264629322488154, - 64'd51461067578504, 64'd617550689667969536, - 64'd25312011692674300, 64'd1252531394179888, - 64'd51374395143744, 64'd604968636770121472, - 64'd25016093697129516, 64'd1240323932807655, - 64'd51271013884936, 64'd592534690332615168, - 64'd24719607558888068, 64'd1228014790252753, - 64'd51151461033318, 64'd580249102199010176, - 64'd24422681573323744, 64'd1215611622371095, - 64'd51016263868528, 64'd568112060983220608, - 64'd24125440374093048, 64'd1203121891965191, - 64'd50865939817425, 64'd556123693884747584, - 64'd23828004995552704, 64'd1190552871739988, - 64'd50700996553661, 64'd544284068472831744, - 64'd23530492934667040, 64'd1177911647241926, - 64'd50521932097946, 64'd532593194439779456, - 64'd23233018212397260, 64'd1165205119780615, - 64'd50329234918947, 64'd521051025323726336, - 64'd22935691434564988, 64'd1152440009332563, - 64'd50123384034768, 64'd509657460201103296, - 64'd22638619852182940, 64'd1139622857426379, - 64'd49904849114947, 64'd498412345349069440, - 64'd22341907421245864, 64'd1126760030008939, - 64'd49674090582925, 64'd487315475878187648, - 64'd22045654861975544, 64'd1113857720291995, - 64'd49431559718931, 64'd476366597335613824, - 64'd21749959717513728, 64'd1100921951578746, - 64'd49177698763229}};
	localparam logic signed[63:0] Fbr[0:3][0:99] = '{
		'{- 64'd209367917907850816, 64'd12940596353402938, 64'd896381733843701, 64'd5773941780322, - 64'd215697698286196160, 64'd12377665357757680, 64'd899926540939321, 64'd6975477820499, - 64'd221744772881992928, 64'd11809873366082668, 64'd902572342792447, 64'd8155642492392, - 64'd227506861175543360, 64'd11237819785294670, 64'd904327652903445, 64'd9313576045912, - 64'd232981981547220352, 64'd10662100720251796, 64'd905201726880791, 64'd10448450412235, - 64'd238168449494480192, 64'd10083308447572872, 64'd905204544538224, 64'd11559469602358, - 64'd243064875588293056, 64'd9502030899551228, 64'd904346791523053, 64'd12645870070256, - 64'd247670163174130496, 64'd8918851158529572, 64'd902639840498836, 64'd13706921040752, - 64'd251983505822829600, 64'd8334346962088413, 64'd900095731905798, 64'd14741924802207, - 64'd256004384536825024, 64'd7749090219385679, 64'd896727154322443, 64'd15750216964190, - 64'd259732564717406848, 64'd7163646538970562, 64'd892547424451934, 64'd16731166680303, - 64'd263168092898817728, 64'd6578574768379709, 64'd887570466756864, 64'd17684176836396, - 64'd266311293255155840, 64'd5994426545808893, 64'd881810792766088, 64'd18608684204390, - 64'd269162763886189760, 64'd5411745864138234, 64'd875283480077328, 64'd19504159562015, - 64'd271723372888330976, 64'd4831068647573912, 64'd868004151079220, 64'd20370107778738, - 64'd273994254217131520, 64'd4252922341153986, 64'd859988951416491, 64'd21206067868235, - 64'd275976803347800640, 64'd3677825513350828, 64'd851254528221888, 64'd22011613007759, - 64'd277672672740341760, 64'd3106287471987255, 64'd841818008138399, 64'd22786350524788, - 64'd279083767116018560, 64'd2538807893668153, 64'd831696975155255, 64'd23529921851380, - 64'd280212238551954656, 64'd1975876466914083, 64'd820909448281046, 64'd24242002446658, - 64'd281060481400761920, 64'd1417972549168047, 64'd809473859077193, 64'd24922301687903, - 64'd281631127042172608, 64'd865564837831255, 64'd797409029074828, 64'd25570562730737, - 64'd281927038473727296, 64'd319111055468575, 64'd784734147098001, 64'd26186562338910, - 64'd281951304747633280, - 64'd220942350690998, 64'd771468746515904, 64'd26770110684226, - 64'd281707235260971136, - 64'd754160494848410, 64'd757632682446620, 64'd27321051117161},
		'{- 64'd209367917907958112, 64'd12940596353398758, 64'd896381733843569, 64'd5773941780326, - 64'd215697698286299968, 64'd12377665357753640, 64'd899926540939193, 64'd6975477820503, - 64'd221744772882093280, 64'd11809873366078768, 64'd902572342792324, 64'd8155642492396, - 64'd227506861175640128, 64'd11237819785290916, 64'd904327652903325, 64'd9313576045915, - 64'd232981981547313472, 64'd10662100720248186, 64'd905201726880675, 64'd10448450412239, - 64'd238168449494569664, 64'd10083308447569412, 64'd905204544538113, 64'd11559469602361, - 64'd243064875588378848, 64'd9502030899547916, 64'd904346791522946, 64'd12645870070259, - 64'd247670163174212544, 64'd8918851158526408, 64'd902639840498734, 64'd13706921040755, - 64'd251983505822907872, 64'd8334346962085402, 64'd900095731905700, 64'd14741924802210, - 64'd256004384536899488, 64'd7749090219382820, 64'd896727154322349, 64'd15750216964192, - 64'd259732564717477504, 64'd7163646538967858, 64'd892547424451845, 64'd16731166680306, - 64'd263168092898884544, 64'd6578574768377158, 64'd887570466756779, 64'd17684176836398, - 64'd266311293255218816, 64'd5994426545806495, 64'd881810792766008, 64'd18608684204392, - 64'd269162763886248896, 64'd5411745864135991, 64'd875283480077252, 64'd19504159562017, - 64'd271723372888386208, 64'd4831068647571824, 64'd868004151079148, 64'd20370107778739, - 64'd273994254217182848, 64'd4252922341152053, 64'd859988951416425, 64'd21206067868237, - 64'd275976803347848064, 64'd3677825513349051, 64'd851254528221826, 64'd22011613007760, - 64'd277672672740385280, 64'd3106287471985634, 64'd841818008138342, 64'd22786350524789, - 64'd279083767116058240, 64'd2538807893666684, 64'd831696975155202, 64'd23529921851382, - 64'd280212238551990528, 64'd1975876466912769, 64'd820909448280998, 64'd24242002446659, - 64'd281060481400793856, 64'd1417972549166887, 64'd809473859077149, 64'd24922301687904, - 64'd281631127042200768, 64'd865564837830247, 64'd797409029074788, 64'd25570562730738, - 64'd281927038473751616, 64'd319111055467717, 64'd784734147097966, 64'd26186562338911, - 64'd281951304747653824, - 64'd220942350691705, 64'd771468746515874, 64'd26770110684226, - 64'd281707235260987936, - 64'd754160494848966, 64'd757632682446594, 64'd27321051117161},
		'{- 64'd208807812964745760, 64'd12908849052433810, 64'd876670745151696, 64'd74765294786063, - 64'd215125675568580832, 64'd12364546145487408, 64'd846574522093956, 64'd73015021252188, - 64'd221174290868974432, 64'd11831835552141554, 64'd817058095947687, 64'd71289534886562, - 64'd226959418591712288, 64'd11310571551516128, 64'd788115257212276, 64'd69588744339475, - 64'd232486745611835648, 64'd10800608470538784, 64'd759739766193057, 64'd67912551711317, - 64'd237761885990934528, 64'd10301800737227882, 64'd731925356245339, 64'd66260852784717, - 64'd242790381040674016, 64'd9814002932348062, 64'd704665736931800, 64'd64633537252140, - 64'd247577699411748000, 64'd9337069839467642, 64'd677954597094628, 64'd63030488938973, - 64'd252129237207467552, 64'd8870856493446672, 64'd651785607843809, 64'd61451586022165, - 64'd256450318121207584, 64'd8415218227384312, 64'd626152425462938, 64'd59896701244465, - 64'd260546193596947328, 64'd7970010718053768, 64'd601048694233914, 64'd58365702124314, - 64'd264422043012156608, 64'd7535090029852914, 64'd576468049181897, 64'd56858451161428, - 64'd268082973882291328, 64'd7110312657298326, 64'd552404118741850, 64'd55374806038149, - 64'd271534022086178720, 64'd6695535566090250, 64'd528850527348025, 64'd53914619816584, - 64'd274780152111582368, 64'd6290616232775662, 64'd505800897947707, 64'd52477741131608, - 64'd277826257320254464, 64'd5895412683036402, 64'd483248854440530, 64'd51064014379769, - 64'd280677160231793856, 64'd5509783528628952, 64'd461188024044683, 64'd49673279904155, - 64'd283337612825642464, 64'd5133588003002269, 64'd439612039591281, 64'd48305374175258, - 64'd285812296860565440, 64'd4766685995619665, 64'd418514541748187, 64'd46960129967909, - 64'd288105824210973600, 64'd4408938085010547, 64'd397889181174568, 64'd45637376534320, - 64'd290222737219459648, 64'd4060205570577469, 64'd377729620607419, 64'd44336939773278, - 64'd292167509064932096, 64'd3720350503183700, 64'd358029536881318, 64'd43058642395570, - 64'd293944544145742976, 64'd3389235714546153, 64'd338782622882642, 64'd41802304085651, - 64'd295558178477218880, 64'd3066724845458330, 64'd319982589439454, 64'd40567741659640, - 64'd297012680103015168, 64'd2752682372867516, 64'd301623167148285, 64'd39354769219676},
		'{- 64'd208807812965074720, 64'd12908849052420436, 64'd876670745151279, 64'd74765294786075, - 64'd215125675568903712, 64'd12364546145474280, 64'd846574522093546, 64'd73015021252200, - 64'd221174290869291296, 64'd11831835552128672, 64'd817058095947284, 64'd71289534886574, - 64'd226959418592023200, 64'd11310571551503488, 64'd788115257211881, 64'd69588744339487, - 64'd232486745612140672, 64'd10800608470526384, 64'd759739766192669, 64'd67912551711329, - 64'd237761885991233696, 64'd10301800737215720, 64'd731925356244959, 64'd66260852784729, - 64'd242790381040967424, 64'd9814002932336134, 64'd704665736931427, 64'd64633537252152, - 64'd247577699412035712, 64'd9337069839455944, 64'd677954597094262, 64'd63030488938984, - 64'd252129237207749632, 64'd8870856493435206, 64'd651785607843450, 64'd61451586022176, - 64'd256450318121484064, 64'd8415218227373072, 64'd626152425462585, 64'd59896701244476, - 64'd260546193597218304, 64'd7970010718042754, 64'd601048694233569, 64'd58365702124324, - 64'd264422043012422080, 64'd7535090029842121, 64'd576468049181558, 64'd56858451161439, - 64'd268082973882551424, 64'd7110312657287754, 64'd552404118741518, 64'd55374806038159, - 64'd271534022086433504, 64'd6695535566079894, 64'd528850527347700, 64'd53914619816594, - 64'd274780152111831872, 64'd6290616232765520, 64'd505800897947388, 64'd52477741131617, - 64'd277826257320498752, 64'd5895412683026470, 64'd483248854440218, 64'd51064014379779, - 64'd280677160232033024, 64'd5509783528619232, 64'd461188024044378, 64'd49673279904164, - 64'd283337612825876544, 64'd5133588002992756, 64'd439612039590981, 64'd48305374175267, - 64'd285812296860794496, 64'd4766685995610355, 64'd418514541747894, 64'd46960129967918, - 64'd288105824211197728, 64'd4408938085001438, 64'd397889181174281, 64'd45637376534328, - 64'd290222737219678848, 64'd4060205570568558, 64'd377729620607138, 64'd44336939773286, - 64'd292167509065146496, 64'd3720350503174987, 64'd358029536881044, 64'd43058642395578, - 64'd293944544145952640, 64'd3389235714537633, 64'd338782622882373, 64'd41802304085659, - 64'd295558178477423808, 64'd3066724845450001, 64'd319982589439191, 64'd40567741659648, - 64'd297012680103215488, 64'd2752682372859375, 64'd301623167148028, 64'd39354769219683}};
	localparam logic signed[63:0] Fbi[0:3][0:99] = '{
		'{64'd256127510662709344, 64'd15852187053065382, - 64'd314423079823242, - 64'd41164091899801, 64'd248129395814423328, 64'd16137135790239808, - 64'd285349582355099, - 64'd40718142853921, 64'd239993514431440960, 64'd16403248028101054, - 64'd256361481670483, - 64'd40238955728992, 64'd231729291000865696, 64'd16650501866890788, - 64'd227485287792818, - 64'd39727393821403, 64'd223346156401711360, 64'd16878893603318750, - 64'd198747079143438, - 64'd39184340614075, 64'd214853538860987136, 64'd17088437510854180, - 64'd170172483044807, - 64'd38610698688936, 64'd206260855023252512, 64'd17279165605622898, - 64'd141786656891765, - 64'd38007388634573, 64'd197577501140738400, 64'd17451127398309160, - 64'd113614270000494, - 64'd37375347950170, 64'd188812844390932416, 64'd17604389632469850, - 64'd85679486144150, - 64'd36715529946819, 64'd179976214328316672, 64'd17739036009676462, - 64'd58005946783340, - 64'd36028902647275, 64'd171076894476740416, 64'd17855166901907766, - 64'd30616754998861, - 64'd35316447685221, 64'd162124114068693760, 64'd17952899051622972, - 64'd3534460133363, - 64'd34579159205100, 64'd153127039937533984, 64'd18032365259951640, 64'd23218956852172, - 64'd33818042763551, 64'd144094768568495984, 64'd18093714063442580, 64'd49622097301960, - 64'd33034114233470, 64'd135036318314095360, 64'd18137109399819340, 64'd75654158064577, - 64'd32228398711708, 64'd125960621779307344, 64'd18162730263194952, 64'd101294943964075, - 64'd31401929431406, 64'd116876518381679152, 64'd18170770349202968, 64'd126524879540126, - 64'd30555746679929, 64'd107792747091301296, 64'd18161437690505888, 64'd151325020055019, - 64'd29690896723379, 64'd98717939355333744, 64'd18134954283145528, 64'd175677061766010, - 64'd28808430738610, 64'd89660612211549136, 64'd18091555704202836, 64'd199563351462307, - 64'd27909403753678, 64'd80629161595120784, 64'd18031490721237340, 64'd222966895266617, - 64'd26994873597632, 64'd71631855842647376, 64'd17955020893978248, 64'd245871366701920, - 64'd26065899860521, 64'd62676829397171616, 64'd17862420168741000, 64'd268261114024824, - 64'd25123542864488, 64'd53772076717708672, 64'd17753974466044040, 64'd290121166827504, - 64'd24168862646791, 64'd44925446396568800, 64'd17629981261901270, 64'd311437241910954, - 64'd23202917955564},
		'{- 64'd256127510662618048, - 64'd15852187053061658, 64'd314423079823345, 64'd41164091899796, - 64'd248129395814329408, - 64'd16137135790235982, 64'd285349582355205, 64'd40718142853917, - 64'd239993514431344512, - 64'd16403248028097132, 64'd256361481670592, 64'd40238955728987, - 64'd231729291000766880, - 64'd16650501866886776, 64'd227485287792931, 64'd39727393821398, - 64'd223346156401610272, - 64'd16878893603314652, 64'd198747079143554, 64'd39184340614070, - 64'd214853538860883936, - 64'd17088437510849998, 64'd170172483044925, 64'd38610698688932, - 64'd206260855023147264, - 64'd17279165605618642, 64'd141786656891886, 64'd38007388634568, - 64'd197577501140631296, - 64'd17451127398304828, 64'd113614270000618, 64'd37375347950165, - 64'd188812844390823520, - 64'd17604389632465452, 64'd85679486144276, 64'd36715529946814, - 64'd179976214328206144, - 64'd17739036009672002, 64'd58005946783468, 64'd36028902647270, - 64'd171076894476628416, - 64'd17855166901903252, 64'd30616754998991, 64'd35316447685216, - 64'd162124114068580352, - 64'd17952899051618404, 64'd3534460133494, 64'd34579159205095, - 64'd153127039937419296, - 64'd18032365259947028, - 64'd23218956852039, 64'd33818042763546, - 64'd144094768568380176, - 64'd18093714063437924, - 64'd49622097301825, 64'd33034114233465, - 64'd135036318313978528, - 64'd18137109399814648, - 64'd75654158064441, 64'd32228398711703, - 64'd125960621779189600, - 64'd18162730263190228, - 64'd101294943963937, 64'd31401929431400, - 64'd116876518381560656, - 64'd18170770349198216, - 64'd126524879539988, 64'd30555746679924, - 64'd107792747091182144, - 64'd18161437690501116, - 64'd151325020054879, 64'd29690896723374, - 64'd98717939355214080, - 64'd18134954283140736, - 64'd175677061765869, 64'd28808430738604, - 64'd89660612211429088, - 64'd18091555704198032, - 64'd199563351462166, 64'd27909403753672, - 64'd80629161595000416, - 64'd18031490721232532, - 64'd222966895266475, 64'd26994873597627, - 64'd71631855842526880, - 64'd17955020893973436, - 64'd245871366701779, 64'd26065899860516, - 64'd62676829397051056, - 64'd17862420168736188, - 64'd268261114024682, 64'd25123542864483, - 64'd53772076717588176, - 64'd17753974466039234, - 64'd290121166827362, 64'd24168862646785, - 64'd44925446396448464, - 64'd17629981261896476, - 64'd311437241910812, 64'd23202917955559},
		'{64'd779901327374593024, 64'd28766736086525376, 64'd1388026451385535, 64'd51147782792348, 64'd765587272939073280, 64'd28489063021489052, 64'd1377710692110832, 64'd51283306989880, 64'd751412666690274560, 64'd28208973279885160, 64'd1367185227349448, 64'd51395528697467, 64'd737378672460398336, 64'd27926644138938352, 64'd1356460265322528, 64'd51485100856128, 64'd723486366557601280, 64'd27642248428922260, 64'd1345545784674669, 64'd51552665436647, 64'd709736739972521728, 64'd27355954600898964, 64'd1334451537574361, 64'd51598853525713, 64'd696130700551027584, 64'd27067926794082408, 64'd1323187052806982, 64'd51624285413561, 64'd682669075133381504, 64'd26778324902811884, 64'd1311761638859439, 64'd51629570683067, 64'd669352611660017792, 64'd26487304643121916, 64'd1300184386995524, 64'd51615308300201, 64'd656181981244139648, 64'd26195017618895720, 64'd1288464174321125, 64'd51582086705768, 64'd643157780211344768, 64'd25901611387589656, 64'd1276609666838425, 64'd51530483908368, 64'd630280532106499840, 64'd25607229525516912, 64'd1264629322488288, 64'd51461067578499, 64'd617550689668085120, 64'd25312011692679012, 64'd1252531394180023, 64'd51374395143739, 64'd604968636770238464, 64'd25016093697134284, 64'd1240323932807792, 64'd51271013884931, 64'd592534690332733568, 64'd24719607558892892, 64'd1228014790252892, 64'd51151461033313, 64'd580249102199129728, 64'd24422681573328616, 64'd1215611622371236, 64'd51016263868523, 64'd568112060983341312, 64'd24125440374097968, 64'd1203121891965334, 64'd50865939817420, 64'd556123693884869504, 64'd23828004995557668, 64'd1190552871740133, 64'd50700996553656, 64'd544284068472954624, 64'd23530492934672044, 64'd1177911647242071, 64'd50521932097940, 64'd532593194439903232, 64'd23233018212402304, 64'd1165205119780762, 64'd50329234918942, 64'd521051025323850944, 64'd22935691434570068, 64'd1152440009332711, 64'd50123384034762, 64'd509657460201228672, 64'd22638619852188048, 64'd1139622857426528, 64'd49904849114941, 64'd498412345349195520, 64'd22341907421251000, 64'd1126760030009089, 64'd49674090582920, 64'd487315475878314432, 64'd22045654861980704, 64'd1113857720292146, 64'd49431559718926, 64'd476366597335741120, 64'd21749959717518912, 64'd1100921951578898, 64'd49177698763224},
		'{- 64'd779901327374501888, - 64'd28766736086521656, - 64'd1388026451385433, - 64'd51147782792353, - 64'd765587272938979456, - 64'd28489063021485228, - 64'd1377710692110726, - 64'd51283306989884, - 64'd751412666690178304, - 64'd28208973279881232, - 64'd1367185227349340, - 64'd51395528697472, - 64'd737378672460299648, - 64'd27926644138934324, - 64'd1356460265322416, - 64'd51485100856132, - 64'd723486366557500416, - 64'd27642248428918144, - 64'd1345545784674554, - 64'd51552665436652, - 64'd709736739972418560, - 64'd27355954600894760, - 64'd1334451537574243, - 64'd51598853525718, - 64'd696130700550922368, - 64'd27067926794078116, - 64'd1323187052806861, - 64'd51624285413566, - 64'd682669075133274368, - 64'd26778324902807512, - 64'd1311761638859315, - 64'd51629570683072, - 64'd669352611659908864, - 64'd26487304643117472, - 64'd1300184386995398, - 64'd51615308300206, - 64'd656181981244028800, - 64'd26195017618891204, - 64'd1288464174320996, - 64'd51582086705773, - 64'd643157780211232128, - 64'd25901611387585068, - 64'd1276609666838294, - 64'd51530483908373, - 64'd630280532106385792, - 64'd25607229525512260, - 64'd1264629322488154, - 64'd51461067578504, - 64'd617550689667969536, - 64'd25312011692674300, - 64'd1252531394179888, - 64'd51374395143744, - 64'd604968636770121472, - 64'd25016093697129516, - 64'd1240323932807655, - 64'd51271013884936, - 64'd592534690332615168, - 64'd24719607558888068, - 64'd1228014790252753, - 64'd51151461033318, - 64'd580249102199010176, - 64'd24422681573323744, - 64'd1215611622371095, - 64'd51016263868528, - 64'd568112060983220608, - 64'd24125440374093048, - 64'd1203121891965191, - 64'd50865939817425, - 64'd556123693884747584, - 64'd23828004995552704, - 64'd1190552871739988, - 64'd50700996553661, - 64'd544284068472831744, - 64'd23530492934667040, - 64'd1177911647241926, - 64'd50521932097946, - 64'd532593194439779456, - 64'd23233018212397260, - 64'd1165205119780615, - 64'd50329234918947, - 64'd521051025323726336, - 64'd22935691434564988, - 64'd1152440009332563, - 64'd50123384034768, - 64'd509657460201103296, - 64'd22638619852182940, - 64'd1139622857426379, - 64'd49904849114947, - 64'd498412345349069440, - 64'd22341907421245864, - 64'd1126760030008939, - 64'd49674090582925, - 64'd487315475878187648, - 64'd22045654861975544, - 64'd1113857720291995, - 64'd49431559718931, - 64'd476366597335613824, - 64'd21749959717513728, - 64'd1100921951578746, - 64'd49177698763229}};
	localparam logic signed[63:0] hf[0:1199] = {64'd2940850143232, - 64'd1165638016, - 64'd1512799744, 64'd1185562, 64'd2939684651008, - 64'd3495991296, - 64'd1510358656, 64'd3554093, 64'd2937354715136, - 64'd5823578112, - 64'd1505480576, 64'd5914922, 64'd2933861908480, - 64'd8146558464, - 64'd1498172544, 64'd8263087, 64'd2929209114624, - 64'd10463097856, - 64'd1488445568, 64'd10593773, 64'd2923400003584, - 64'd12771369984, - 64'd1476313728, 64'd12902316, 64'd2916439293952, - 64'd15069559808, - 64'd1461794304, 64'd15184202, 64'd2908332490752, - 64'd17355862016, - 64'd1444908160, 64'd17435072, 64'd2899085885440, - 64'd19628486656, - 64'd1425678720, 64'd19650720, 64'd2888706555904, - 64'd21885661184, - 64'd1404132736, 64'd21827094, 64'd2877203152896, - 64'd24125630464, - 64'd1380300032, 64'd23960296, 64'd2864584065024, - 64'd26346659840, - 64'd1354212864, 64'd26046590, 64'd2850859778048, - 64'd28547035136, - 64'd1325906688, 64'd28082390, 64'd2836040777728, - 64'd30725066752, - 64'd1295419264, 64'd30064270, 64'd2820138860544, - 64'd32879091712, - 64'd1262791040, 64'd31988960, 64'd2803166085120, - 64'd35007475712, - 64'd1228064896, 64'd33853348, 64'd2785135820800, - 64'd37108604928, - 64'd1191286400, 64'd35654480, 64'd2766062223360, - 64'd39180910592, - 64'd1152503040, 64'd37389556, 64'd2745959972864, - 64'd41222840320, - 64'd1111764480, 64'd39055932, 64'd2724844797952, - 64'd43232890880, - 64'd1069122880, 64'd40651128, 64'd2702732689408, - 64'd45209579520, - 64'd1024631936, 64'd42172808, 64'd2679640948736, - 64'd47151468544, - 64'd978347520, 64'd43618800, 64'd2655587139584, - 64'd49057153024, - 64'd930327232, 64'd44987076, 64'd2630589874176, - 64'd50925277184, - 64'd880630464, 64'd46275772, 64'd2604668289024, - 64'd52754509824, - 64'd829318080, 64'd47483168, 64'd2577842307072, - 64'd54543568896, - 64'd776452544, 64'd48607692, 64'd2550131851264, - 64'd56291221504, - 64'd722097728, 64'd49647932, 64'd2521558155264, - 64'd57996267520, - 64'd666318784, 64'd50602608, 64'd2492142714880, - 64'd59657555968, - 64'd609182208, 64'd51470604, 64'd2461908074496, - 64'd61273976832, - 64'd550755456, 64'd52250928, 64'd2430876516352, - 64'd62844473344, - 64'd491107104, 64'd52942748, 64'd2399071371264, - 64'd64368029696, - 64'd430306720, 64'd53545364, 64'd2366516494336, - 64'd65843679232, - 64'd368424576, 64'd54058212, 64'd2333235740672, - 64'd67270504448, - 64'd305531808, 64'd54480872, 64'd2299254276096, - 64'd68647636992, - 64'd241700112, 64'd54813048, 64'd2264596480000, - 64'd69974253568, - 64'd177001840, 64'd55054588, 64'd2229288566784, - 64'd71249592320, - 64'd111509720, 64'd55205460, 64'd2193355702272, - 64'd72472920064, - 64'd45296908, 64'd55265764, 64'd2156824363008, - 64'd73643573248, 64'd21563162, 64'd55235720, 64'd2119720894464, - 64'd74760937472, 64'd88996872, 64'd55115676, 64'd2082072297472, - 64'd75824447488, 64'd156930480, 64'd54906092, 64'd2043905572864, - 64'd76833570816, 64'd225290224, 64'd54607548, 64'd2005247983616, - 64'd77787865088, 64'd294002400, 64'd54220744, 64'd1966126923776, - 64'd78686896128, 64'd362993504, 64'd53746476, 64'd1926570311680, - 64'd79530311680, 64'd432190112, 64'd53185660, 64'd1886605934592, - 64'd80317808640, 64'd501519296, 64'd52539316, 64'd1846261841920, - 64'd81049116672, 64'd570908416, 64'd51808560, 64'd1805566214144, - 64'd81724030976, 64'd640285248, 64'd50994608, 64'd1764547231744, - 64'd82342395904, 64'd709578176, 64'd50098780, 64'd1723233206272, - 64'd82904104960, 64'd778716288, 64'd49122472, 64'd1681652580352, - 64'd83409100800, 64'd847629120, 64'd48067184, 64'd1639833665536, - 64'd83857383424, 64'd916247232, 64'd46934500, 64'd1597804642304, - 64'd84249001984, 64'd984501824, 64'd45726076, 64'd1555594084352, - 64'd84584038400, 64'd1052325120, 64'd44443660, 64'd1513230041088, - 64'd84862640128, 64'd1119650176, 64'd43089068, 64'd1470740824064, - 64'd85084995584, 64'd1186411136, 64'd41664192, 64'd1428154351616, - 64'd85251350528, 64'd1252543232, 64'd40170992, 64'd1385498673152, - 64'd85361983488, 64'd1317982720, 64'd38611496, 64'd1342801575936, - 64'd85417230336, 64'd1382667392, 64'd36987788, 64'd1300090585088, - 64'd85417467904, 64'd1446536064, 64'd35302024, 64'd1257393225728, - 64'd85363122176, 64'd1509528704, 64'd33556404, 64'd1214736498688, - 64'd85254660096, 64'd1571586816, 64'd31753180, 64'd1172147535872, - 64'd85092589568, 64'd1632653312, 64'd29894662, 64'd1129652813824, - 64'd84877467648, 64'd1692672640, 64'd27983200, 64'd1087278809088, - 64'd84609875968, 64'd1751590528, 64'd26021184, 64'd1045051539456, - 64'd84290469888, 64'd1809354496, 64'd24011048, 64'd1002996826112, - 64'd83919912960, 64'd1865913472, 64'd21955256, 64'd961140031488, - 64'd83498917888, 64'd1921217920, 64'd19856308, 64'd919506190336, - 64'd83028238336, 64'd1975220352, 64'd17716730, 64'd878119944192, - 64'd82508668928, 64'd2027874432, 64'd15539076, 64'd837005541376, - 64'd81941028864, 64'd2079135872, 64'd13325920, 64'd796186771456, - 64'd81326186496, 64'd2128962048, 64'd11079857, 64'd755687096320, - 64'd80665018368, 64'd2177312256, 64'd8803495, 64'd715529322496, - 64'd79958450176, 64'd2224147456, 64'd6499455, 64'd675736059904, - 64'd79207456768, 64'd2269430272, 64'd4170370, 64'd636329132032, - 64'd78413004800, 64'd2313125632, 64'd1818876, 64'd597330100224, - 64'd77576118272, 64'd2355199744, - 64'd552387, 64'd558759936000, - 64'd76697837568, 64'd2395620864, - 64'd2940777, 64'd520638988288, - 64'd75779235840, 64'd2434359808, - 64'd5343657, 64'd482987212800, - 64'd74821394432, 64'd2471388160, - 64'd7758395, 64'd445823942656, - 64'd73825452032, 64'd2506680320, - 64'd10182368, 64'd409167921152, - 64'd72792530944, 64'd2540212224, - 64'd12612964, 64'd373037367296, - 64'd71723802624, 64'd2571961600, - 64'd15047585, 64'd337449910272, - 64'd70620454912, 64'd2601908224, - 64'd17483650, 64'd302422491136, - 64'd69483675648, 64'd2630034432, - 64'd19918600, 64'd267971592192, - 64'd68314685440, 64'd2656323072, - 64'd22349896, 64'd234112974848, - 64'd67114729472, 64'd2680760576, - 64'd24775022, 64'd200861810688, - 64'd65885052928, 64'd2703333888, - 64'd27191490, 64'd168232665088, - 64'd64626917376, 64'd2724032768, - 64'd29596848, 64'd136239431680, - 64'd63341600768, 64'd2742848256, - 64'd31988666, 64'd104895381504, - 64'd62030393344, 64'd2759773952, - 64'd34364556, 64'd74213138432, - 64'd60694589440, 64'd2774804736, - 64'd36722164, 64'd44204675072, - 64'd59335491584, 64'd2787937536, - 64'd39059168, 64'd14881307648, - 64'd57954418688, 64'd2799171328, - 64'd41373300, - 64'd13746302976, - 64'd56552689664, 64'd2808506880, - 64'd43662328, - 64'd41668161536, - 64'd55131627520, 64'd2815946496, - 64'd45924056, - 64'd68874928128, - 64'd53692555264, 64'd2821494528, - 64'd48156352, - 64'd95357935616, - 64'd52236808192, 64'd2825156864, - 64'd50357112, - 64'd121109176320, - 64'd50765713408, 64'd2826941696, - 64'd52524304, - 64'd146121310208, - 64'd49280606208, 64'd2826857984, - 64'd54655932, - 64'd170387668992, - 64'd47782809600, 64'd2824917504, - 64'd56750052, - 64'd193902231552, - 64'd46273650688, 64'd2821132800, - 64'd58804788, - 64'd216659656704, - 64'd44754456576, 64'd2815518464, - 64'd60818304, - 64'd238655242240, - 64'd43226542080, 64'd2808090624, - 64'd62788840, - 64'd259884957696, - 64'd41691217920, 64'd2798866944, - 64'd64714672, - 64'd280345444352, - 64'd40149786624, 64'd2787866880, - 64'd66594152, - 64'd300033933312, - 64'd38603550720, 64'd2775110912, - 64'd68425696, - 64'd318948409344, - 64'd37053788160, 64'd2760621312, - 64'd70207760, - 64'd337087365120, - 64'd35501780992, 64'd2744421888, - 64'd71938888, - 64'd354450014208, - 64'd33948788736, 64'd2726537728, - 64'd73617664, - 64'd371036192768, - 64'd32396066816, 64'd2706995200, - 64'd75242768, - 64'd386846326784, - 64'd30844850176, 64'd2685821696, - 64'd76812912, - 64'd401881497600, - 64'd29296365568, 64'd2663046912, - 64'd78326888, - 64'd416143343616, - 64'd27751819264, 64'd2638700544, - 64'd79783560, - 64'd429634158592, - 64'd26212401152, 64'd2612814336, - 64'd81181848, - 64'd442356793344, - 64'd24679286784, 64'd2585420544, - 64'd82520744, - 64'd454314688512, - 64'd23153633280, 64'd2556553472, - 64'd83799312, - 64'd465511874560, - 64'd21636573184, 64'd2526247424, - 64'd85016672, - 64'd475952873472, - 64'd20129226752, 64'd2494538240, - 64'd86172024, - 64'd485642895360, - 64'd18632689664, 64'd2461462784, - 64'd87264632, - 64'd494587543552, - 64'd17148034048, 64'd2427058944, - 64'd88293824, - 64'd502793076736, - 64'd15676313600, 64'd2391365376, - 64'd89259000, - 64'd510266212352, - 64'd14218556416, 64'd2354420992, - 64'd90159632, - 64'd517014126592, - 64'd12775770112, 64'd2316266496, - 64'd90995240, - 64'd523044618240, - 64'd11348933632, 64'd2276942592, - 64'd91765448, - 64'd528365879296, - 64'd9939003392, 64'd2236491264, - 64'd92469904, - 64'd532986593280, - 64'd8546911744, 64'd2194954752, - 64'd93108368, - 64'd536915935232, - 64'd7173561856, 64'd2152375552, - 64'd93680616, - 64'd540163440640, - 64'd5819831808, 64'd2108797824, - 64'd94186544, - 64'd542739169280, - 64'd4486573056, 64'd2064265216, - 64'd94626064, - 64'd544653541376, - 64'd3174608640, 64'd2018822272, - 64'd94999192, - 64'd545917468672, - 64'd1884733568, 64'd1972513664, - 64'd95305976, - 64'd546542092288, - 64'd617714624, 64'd1925384960, - 64'd95546560, - 64'd546539110400, 64'd625710208, 64'd1877481600, - 64'd95721120, - 64'd545920450560, 64'd1844832128, 64'd1828849408, - 64'd95829912, - 64'd544698433536, 64'd3038971904, 64'd1779534464, - 64'd95873240, - 64'd542885740544, 64'd4207480064, 64'd1729583104, - 64'd95851488, - 64'd540495314944, 64'd5349736960, 64'd1679041664, - 64'd95765088, - 64'd537540460544, 64'd6465153536, 64'd1627956480, - 64'd95614512, - 64'd534034743296, 64'd7553170944, 64'd1576374400, - 64'd95400320, - 64'd529991958528, 64'd8613261312, 64'd1524341760, - 64'd95123112, - 64'd525426229248, 64'd9644926976, 64'd1471905024, - 64'd94783544, - 64'd520351842304, 64'd10647700480, 64'd1419110784, - 64'd94382320, - 64'd514783412224, 64'd11621147648, 64'd1366005120, - 64'd93920200, - 64'd508735651840, 64'd12564862976, 64'd1312634368, - 64'd93398000, - 64'd502223568896, 64'd13478472704, 64'd1259044096, - 64'd92816584, - 64'd495262269440, 64'd14361633792, 64'd1205280256, - 64'd92176856, - 64'd487867056128, 64'd15214034944, 64'd1151388032, - 64'd91479784, - 64'd480053395456, 64'd16035394560, 64'd1097412480, - 64'd90726352, - 64'd471836884992, 64'd16825462784, 64'd1043398272, - 64'd89917624, - 64'd463233187840, 64'd17584019456, 64'd989389632, - 64'd89054672, - 64'd454258130944, 64'd18310875136, 64'd935430336, - 64'd88138632, - 64'd444927606784, 64'd19005870080, 64'd881563648, - 64'd87170672, - 64'd435257606144, 64'd19668875264, 64'd827832448, - 64'd86152000, - 64'd425264087040, 64'd20299794432, 64'd774278848, - 64'd85083856, - 64'd414963171328, 64'd20898553856, 64'd720944576, - 64'd83967520, - 64'd404370915328, 64'd21465116672, 64'd667870656, - 64'd82804296, - 64'd393503408128, 64'd21999468544, 64'd615097408, - 64'd81595528, - 64'd382376804352, 64'd22501629952, 64'd562664512, - 64'd80342592, - 64'd371007160320, 64'd22971641856, 64'd510611008, - 64'd79046888, - 64'd359410499584, 64'd23409582080, 64'd458975104, - 64'd77709832, - 64'd347602878464, 64'd23815548928, 64'd407794272, - 64'd76332888, - 64'd335600254976, 64'd24189671424, 64'd357105184, - 64'd74917520, - 64'd323418488832, 64'd24532105216, 64'd306943680, - 64'd73465224, - 64'd311073406976, 64'd24843030528, 64'd257344752, - 64'd71977528, - 64'd298580672512, 64'd25122652160, 64'd208342576, - 64'd70455960, - 64'd285955948544, 64'd25371203584, 64'd159970368, - 64'd68902072, - 64'd273214619648, 64'd25588940800, 64'd112260464, - 64'd67317424, - 64'd260372086784, 64'd25776146432, 64'd65244268, - 64'd65703596, - 64'd247443505152, 64'd25933123584, 64'd18952236, - 64'd64062188, - 64'd234443948032, 64'd26060197888, - 64'd26586158, - 64'd62394792, - 64'd221388242944, 64'd26157721600, - 64'd71342424, - 64'd60703024, - 64'd208291086336, 64'd26226067456, - 64'd115289064, - 64'd58988492, - 64'd195166978048, 64'd26265624576, - 64'd158399616, - 64'd57252828, - 64'd182030188544, 64'd26276810752, - 64'd200648608, - 64'd55497648, - 64'd168894824448, 64'd26260058112, - 64'd242011664, - 64'd53724580, - 64'd155774713856, 64'd26215821312, - 64'd282465440, - 64'd51935256, - 64'd142683504640, 64'd26144571392, - 64'd321987616, - 64'd50131300, - 64'd129634557952, 64'd26046797824, - 64'd360556992, - 64'd48314332, - 64'd116641038336, 64'd25923008512, - 64'd398153440, - 64'd46485976, - 64'd103715799040, 64'd25773729792, - 64'd434757920, - 64'd44647844, - 64'd90871463936, 64'd25599500288, - 64'd470352448, - 64'd42801540, - 64'd78120370176, 64'd25400875008, - 64'd504920192, - 64'd40948668, - 64'd65474560000, 64'd25178427392, - 64'd538445376, - 64'd39090812, - 64'd52945813504, 64'd24932741120, - 64'd570913344, - 64'd37229548, - 64'd40545595392, 64'd24664412160, - 64'd602310528, - 64'd35366440, - 64'd28285073408, 64'd24374052864, - 64'd632624512, - 64'd33503040, - 64'd16175110144, 64'd24062283776, - 64'd661843904, - 64'd31640880, - 64'd4226252032, 64'd23729739776, - 64'd689958528, - 64'd29781480, 64'd7551273984, 64'd23377063936, - 64'd716959168, - 64'd27926338, 64'd19147565056, 64'd23004909568, - 64'd742837760, - 64'd26076936, 64'd30553047040, 64'd22613938176, - 64'd767587328, - 64'd24234734, 64'd41758478336, 64'd22204823552, - 64'd791202048, - 64'd22401170, 64'd52754960384, 64'd21778241536, - 64'd813677120, - 64'd20577660, 64'd63533924352, 64'd21334876160, - 64'd835008704, - 64'd18765600, 64'd74087153664, 64'd20875419648, - 64'd855194176, - 64'd16966354, 64'd84406779904, 64'd20400570368, - 64'd874231936, - 64'd15181266, 64'd94485274624, 64'd19911026688, - 64'd892121408, - 64'd13411651, 64'd104315469824, 64'd19407495168, - 64'd908862912, - 64'd11658797, 64'd113890557952, 64'd18890684416, - 64'd924457984, - 64'd9923964, 64'd123204067328, 64'd18361305088, - 64'd938909120, - 64'd8208380, 64'd132249886720, 64'd17820069888, - 64'd952219648, - 64'd6513247, 64'd141022281728, 64'd17267693568, - 64'd964394112, - 64'd4839731, 64'd149515845632, 64'd16704888832, - 64'd975437760, - 64'd3188970, 64'd157725540352, 64'd16132372480, - 64'd985357056, - 64'd1562069, 64'd165646712832, 64'd15550857216, - 64'd994159104, 64'd39902, 64'd173275021312, 64'd14961054720, - 64'd1001852224, 64'd1615906, 64'd180606500864, 64'd14363675648, - 64'd1008445312, 64'd3164939, 64'd187637547008, 64'd13759428608, - 64'd1013948352, 64'd4686034, 64'd194364899328, 64'd13149016064, - 64'd1018372160, 64'd6178258, 64'd200785657856, 64'd12533139456, - 64'd1021728256, 64'd7640716, 64'd206897250304, 64'd11912493056, - 64'd1024029120, 64'd9072546, 64'd212697464832, 64'd11287769088, - 64'd1025287936, 64'd10472925, 64'd218184450048, 64'd10659650560, - 64'd1025518720, 64'd11841068, 64'd223356665856, 64'd10028817408, - 64'd1024736192, 64'd13176226, 64'd228212932608, 64'd9395940352, - 64'd1022955776, 64'd14477687, 64'd232752381952, 64'd8761683968, - 64'd1020193664, 64'd15744778, 64'd236974489600, 64'd8126705152, - 64'd1016466752, 64'd16976866, 64'd240879075328, 64'd7491652096, - 64'd1011792384, 64'd18173352, 64'd244466237440, 64'd6857163264, - 64'd1006188864, 64'd19333680, 64'd247736434688, 64'd6223868928, - 64'd999674816, 64'd20457330, 64'd250690404352, 64'd5592388608, - 64'd992269568, 64'd21543820, 64'd253329227776, 64'd4963332608, - 64'd983993088, 64'd22592710, 64'd255654248448, 64'd4337299456, - 64'd974865728, 64'd23603594, 64'd257667121152, 64'd3714877184, - 64'd964908416, 64'd24576108, 64'd259369828352, 64'd3096642048, - 64'd954142592, 64'd25509924, 64'd260764565504, 64'd2483158272, - 64'd942590080, 64'd26404754, 64'd261853855744, 64'd1874978048, - 64'd930273216, 64'd27260348, 64'd262640517120, 64'd1272640384, - 64'd917214656, 64'd28076494, 64'd263127564288, 64'd676671872, - 64'd903437632, 64'd28853018, 64'd263318339584, 64'd87585424, - 64'd888965376, 64'd29589780, 64'd263216381952, - 64'd494119680, - 64'd873821888, 64'd30286680, 64'd262825525248, - 64'd1067958016, - 64'd858031040, 64'd30943656, 64'd262149816320, - 64'd1633458304, - 64'd841617344, 64'd31560682, 64'd261193531392, - 64'd2190163968, - 64'd824605312, 64'd32137764, 64'd259961192448, - 64'd2737633280, - 64'd807019840, 64'd32674948, 64'd258457501696, - 64'd3275438592, - 64'd788885952, 64'd33172316, 64'd256687423488, - 64'd3803168512, - 64'd770228800, 64'd33629976, 64'd254656086016, - 64'd4320425984, - 64'd751073856, 64'd34048084, 64'd252368814080, - 64'd4826830848, - 64'd731446464, 64'd34426820, 64'd249831129088, - 64'd5322016768, - 64'd711372288, 64'd34766396, 64'd247048716288, - 64'd5805634560, - 64'd690876992, 64'd35067064, 64'd244027473920, - 64'd6277350912, - 64'd669986240, 64'd35329100, 64'd240773414912, - 64'd6736847872, - 64'd648725760, 64'd35552820, 64'd237292716032, - 64'd7183823872, - 64'd627121344, 64'd35738560, 64'd233591717888, - 64'd7617994240, - 64'd605198656, 64'd35886692, 64'd229676892160, - 64'd8039089664, - 64'd582983360, 64'd35997620, 64'd225554857984, - 64'd8446857728, - 64'd560501120, 64'd36071772, 64'd221232300032, - 64'd8841062400, - 64'd537777344, 64'd36109608, 64'd216716083200, - 64'd9221482496, - 64'd514837408, 64'd36111604, 64'd212013154304, - 64'd9587915776, - 64'd491706656, 64'd36078280, 64'd207130525696, - 64'd9940173824, - 64'd468410144, 64'd36010168, 64'd202075373568, - 64'd10278087680, - 64'd444972768, 64'd35907824, 64'd196854857728, - 64'd10601500672, - 64'd421419264, 64'd35771840, 64'd191476301824, - 64'd10910274560, - 64'd397774112, 64'd35602824, 64'd185947045888, - 64'd11204287488, - 64'd374061536, 64'd35401396, 64'd180274495488, - 64'd11483432960, - 64'd350305568, 64'd35168220, 64'd174466105344, - 64'd11747620864, - 64'd326529888, 64'd34903956, 64'd168529379328, - 64'd11996775424, - 64'd302757952, 64'd34609308, 64'd162471854080, - 64'd12230838272, - 64'd279012800, 64'd34284976, 64'd156301066240, - 64'd12449766400, - 64'd255317248, 64'd33931692, 64'd150024601600, - 64'd12653530112, - 64'd231693680, 64'd33550202, 64'd143650062336, - 64'd12842118144, - 64'd208164128, 64'd33141266, 64'd137185017856, - 64'd13015530496, - 64'd184750272, 64'd32705664, 64'd130637062144, - 64'd13173785600, - 64'd161473392, 64'd32244184, 64'd124013756416, - 64'd13316914176, - 64'd138354304, 64'd31757632, 64'd117322661888, - 64'd13444962304, - 64'd115413440, 64'd31246826, 64'd110571298816, - 64'd13557988352, - 64'd92670792, 64'd30712592, 64'd103767162880, - 64'd13656068096, - 64'd70145880, 64'd30155772, 64'd96917708800, - 64'd13739287552, - 64'd47857776, 64'd29577214, 64'd90030333952, - 64'd13807748096, - 64'd25825048, 64'd28977778, 64'd83112402944, - 64'd13861564416, - 64'd4065793, 64'd28358328, 64'd76171190272, - 64'd13900861440, 64'd17402396, 64'd27719738, 64'd69213937664, - 64'd13925779456, 64'd38562440, 64'd27062890, 64'd62247784448, - 64'd13936468992, 64'd59397776, 64'd26388666, 64'd55279808512, - 64'd13933095936, 64'd79892376, 64'd25697958, 64'd48317001728, - 64'd13915833344, 64'd100030752, 64'd24991658, 64'd41366261760, - 64'd13884868608, 64'd119797944, 64'd24270660, 64'd34434383872, - 64'd13840399360, 64'd139179568, 64'd23535864, 64'd27528077312, - 64'd13782632448, 64'd158161776, 64'd22788168, 64'd20653932544, - 64'd13711788032, 64'd176731296, 64'd22028472, 64'd13818431488, - 64'd13628093440, 64'd194875424, 64'd21257672, 64'd7027940352, - 64'd13531788288, 64'd212582048, 64'd20476664, 64'd288703872, - 64'd13423118336, 64'd229839616, 64'd19686344, - 64'd6393159680, - 64'd13302340608, 64'd246637136, 64'd18887604, - 64'd13011662848, - 64'd13169720320, 64'd262964256, 64'd18081328, - 64'd19560951808, - 64'd13025530880, 64'd278811168, 64'd17268400, - 64'd26035312640, - 64'd12870052864, 64'd294168672, 64'd16449699, - 64'd32429170688, - 64'd12703575040, 64'd309028160, 64'd15626094, - 64'd38737104896, - 64'd12526392320, 64'd323381600, 64'd14798449, - 64'd44953829376, - 64'd12338807808, 64'd337221536, 64'd13967621, - 64'd51074228224, - 64'd12141129728, 64'd350541152, 64'd13134456, - 64'd57093328896, - 64'd11933672448, 64'd363334208, 64'd12299796, - 64'd63006322688, - 64'd11716757504, 64'd375595008, 64'd11464468, - 64'd68808564736, - 64'd11490709504, 64'd387318496, 64'd10629291, - 64'd74495565824, - 64'd11255858176, 64'd398500160, 64'd9795073, - 64'd80063012864, - 64'd11012540416, 64'd409136096, 64'd8962611, - 64'd85506752512, - 64'd10761092096, 64'd419222944, 64'd8132689, - 64'd90822803456, - 64'd10501858304, 64'd428757984, 64'd7306078, - 64'd96007372800, - 64'd10235184128, 64'd437738944, 64'd6483536};
	localparam logic signed[63:0] hb[0:1199] = {64'd2940850143232, 64'd1165638016, - 64'd1512799744, - 64'd1185562, 64'd2939684651008, 64'd3495991296, - 64'd1510358656, - 64'd3554093, 64'd2937354715136, 64'd5823578112, - 64'd1505480576, - 64'd5914922, 64'd2933861908480, 64'd8146558464, - 64'd1498172544, - 64'd8263087, 64'd2929209114624, 64'd10463097856, - 64'd1488445568, - 64'd10593773, 64'd2923400003584, 64'd12771369984, - 64'd1476313728, - 64'd12902316, 64'd2916439293952, 64'd15069559808, - 64'd1461794304, - 64'd15184202, 64'd2908332490752, 64'd17355862016, - 64'd1444908160, - 64'd17435072, 64'd2899085885440, 64'd19628486656, - 64'd1425678720, - 64'd19650720, 64'd2888706555904, 64'd21885661184, - 64'd1404132736, - 64'd21827094, 64'd2877203152896, 64'd24125630464, - 64'd1380300032, - 64'd23960296, 64'd2864584065024, 64'd26346659840, - 64'd1354212864, - 64'd26046590, 64'd2850859778048, 64'd28547035136, - 64'd1325906688, - 64'd28082390, 64'd2836040777728, 64'd30725066752, - 64'd1295419264, - 64'd30064270, 64'd2820138860544, 64'd32879091712, - 64'd1262791040, - 64'd31988960, 64'd2803166085120, 64'd35007475712, - 64'd1228064896, - 64'd33853348, 64'd2785135820800, 64'd37108604928, - 64'd1191286400, - 64'd35654480, 64'd2766062223360, 64'd39180910592, - 64'd1152503040, - 64'd37389556, 64'd2745959972864, 64'd41222840320, - 64'd1111764480, - 64'd39055932, 64'd2724844797952, 64'd43232890880, - 64'd1069122880, - 64'd40651128, 64'd2702732689408, 64'd45209579520, - 64'd1024631936, - 64'd42172808, 64'd2679640948736, 64'd47151468544, - 64'd978347520, - 64'd43618800, 64'd2655587139584, 64'd49057153024, - 64'd930327232, - 64'd44987076, 64'd2630589874176, 64'd50925277184, - 64'd880630464, - 64'd46275772, 64'd2604668289024, 64'd52754509824, - 64'd829318080, - 64'd47483168, 64'd2577842307072, 64'd54543568896, - 64'd776452544, - 64'd48607692, 64'd2550131851264, 64'd56291221504, - 64'd722097728, - 64'd49647932, 64'd2521558155264, 64'd57996267520, - 64'd666318784, - 64'd50602608, 64'd2492142714880, 64'd59657555968, - 64'd609182208, - 64'd51470604, 64'd2461908074496, 64'd61273976832, - 64'd550755456, - 64'd52250928, 64'd2430876516352, 64'd62844473344, - 64'd491107104, - 64'd52942748, 64'd2399071371264, 64'd64368029696, - 64'd430306720, - 64'd53545364, 64'd2366516494336, 64'd65843679232, - 64'd368424576, - 64'd54058212, 64'd2333235740672, 64'd67270504448, - 64'd305531808, - 64'd54480872, 64'd2299254276096, 64'd68647636992, - 64'd241700112, - 64'd54813048, 64'd2264596480000, 64'd69974253568, - 64'd177001840, - 64'd55054588, 64'd2229288566784, 64'd71249592320, - 64'd111509720, - 64'd55205460, 64'd2193355702272, 64'd72472920064, - 64'd45296908, - 64'd55265764, 64'd2156824363008, 64'd73643573248, 64'd21563162, - 64'd55235720, 64'd2119720894464, 64'd74760937472, 64'd88996872, - 64'd55115676, 64'd2082072297472, 64'd75824447488, 64'd156930480, - 64'd54906092, 64'd2043905572864, 64'd76833570816, 64'd225290224, - 64'd54607548, 64'd2005247983616, 64'd77787865088, 64'd294002400, - 64'd54220744, 64'd1966126923776, 64'd78686896128, 64'd362993504, - 64'd53746476, 64'd1926570311680, 64'd79530311680, 64'd432190112, - 64'd53185660, 64'd1886605934592, 64'd80317808640, 64'd501519296, - 64'd52539316, 64'd1846261841920, 64'd81049116672, 64'd570908416, - 64'd51808560, 64'd1805566214144, 64'd81724030976, 64'd640285248, - 64'd50994608, 64'd1764547231744, 64'd82342395904, 64'd709578176, - 64'd50098780, 64'd1723233206272, 64'd82904104960, 64'd778716288, - 64'd49122472, 64'd1681652580352, 64'd83409100800, 64'd847629120, - 64'd48067184, 64'd1639833665536, 64'd83857383424, 64'd916247232, - 64'd46934500, 64'd1597804642304, 64'd84249001984, 64'd984501824, - 64'd45726076, 64'd1555594084352, 64'd84584038400, 64'd1052325120, - 64'd44443660, 64'd1513230041088, 64'd84862640128, 64'd1119650176, - 64'd43089068, 64'd1470740824064, 64'd85084995584, 64'd1186411136, - 64'd41664192, 64'd1428154351616, 64'd85251350528, 64'd1252543232, - 64'd40170992, 64'd1385498673152, 64'd85361983488, 64'd1317982720, - 64'd38611496, 64'd1342801575936, 64'd85417230336, 64'd1382667392, - 64'd36987788, 64'd1300090585088, 64'd85417467904, 64'd1446536064, - 64'd35302024, 64'd1257393225728, 64'd85363122176, 64'd1509528704, - 64'd33556404, 64'd1214736498688, 64'd85254660096, 64'd1571586816, - 64'd31753180, 64'd1172147535872, 64'd85092589568, 64'd1632653312, - 64'd29894662, 64'd1129652813824, 64'd84877467648, 64'd1692672640, - 64'd27983200, 64'd1087278809088, 64'd84609875968, 64'd1751590528, - 64'd26021184, 64'd1045051539456, 64'd84290469888, 64'd1809354496, - 64'd24011048, 64'd1002996826112, 64'd83919912960, 64'd1865913472, - 64'd21955256, 64'd961140031488, 64'd83498917888, 64'd1921217920, - 64'd19856308, 64'd919506190336, 64'd83028238336, 64'd1975220352, - 64'd17716730, 64'd878119944192, 64'd82508668928, 64'd2027874432, - 64'd15539076, 64'd837005541376, 64'd81941028864, 64'd2079135872, - 64'd13325920, 64'd796186771456, 64'd81326186496, 64'd2128962048, - 64'd11079857, 64'd755687096320, 64'd80665018368, 64'd2177312256, - 64'd8803495, 64'd715529322496, 64'd79958450176, 64'd2224147456, - 64'd6499455, 64'd675736059904, 64'd79207456768, 64'd2269430272, - 64'd4170370, 64'd636329132032, 64'd78413004800, 64'd2313125632, - 64'd1818876, 64'd597330100224, 64'd77576118272, 64'd2355199744, 64'd552387, 64'd558759936000, 64'd76697837568, 64'd2395620864, 64'd2940777, 64'd520638988288, 64'd75779235840, 64'd2434359808, 64'd5343657, 64'd482987212800, 64'd74821394432, 64'd2471388160, 64'd7758395, 64'd445823942656, 64'd73825452032, 64'd2506680320, 64'd10182368, 64'd409167921152, 64'd72792530944, 64'd2540212224, 64'd12612964, 64'd373037367296, 64'd71723802624, 64'd2571961600, 64'd15047585, 64'd337449910272, 64'd70620454912, 64'd2601908224, 64'd17483650, 64'd302422491136, 64'd69483675648, 64'd2630034432, 64'd19918600, 64'd267971592192, 64'd68314685440, 64'd2656323072, 64'd22349896, 64'd234112974848, 64'd67114729472, 64'd2680760576, 64'd24775022, 64'd200861810688, 64'd65885052928, 64'd2703333888, 64'd27191490, 64'd168232665088, 64'd64626917376, 64'd2724032768, 64'd29596848, 64'd136239431680, 64'd63341600768, 64'd2742848256, 64'd31988666, 64'd104895381504, 64'd62030393344, 64'd2759773952, 64'd34364556, 64'd74213138432, 64'd60694589440, 64'd2774804736, 64'd36722164, 64'd44204675072, 64'd59335491584, 64'd2787937536, 64'd39059168, 64'd14881307648, 64'd57954418688, 64'd2799171328, 64'd41373300, - 64'd13746302976, 64'd56552689664, 64'd2808506880, 64'd43662328, - 64'd41668161536, 64'd55131627520, 64'd2815946496, 64'd45924056, - 64'd68874928128, 64'd53692555264, 64'd2821494528, 64'd48156352, - 64'd95357935616, 64'd52236808192, 64'd2825156864, 64'd50357112, - 64'd121109176320, 64'd50765713408, 64'd2826941696, 64'd52524304, - 64'd146121310208, 64'd49280606208, 64'd2826857984, 64'd54655932, - 64'd170387668992, 64'd47782809600, 64'd2824917504, 64'd56750052, - 64'd193902231552, 64'd46273650688, 64'd2821132800, 64'd58804788, - 64'd216659656704, 64'd44754456576, 64'd2815518464, 64'd60818304, - 64'd238655242240, 64'd43226542080, 64'd2808090624, 64'd62788840, - 64'd259884957696, 64'd41691217920, 64'd2798866944, 64'd64714672, - 64'd280345444352, 64'd40149786624, 64'd2787866880, 64'd66594152, - 64'd300033933312, 64'd38603550720, 64'd2775110912, 64'd68425696, - 64'd318948409344, 64'd37053788160, 64'd2760621312, 64'd70207760, - 64'd337087365120, 64'd35501780992, 64'd2744421888, 64'd71938888, - 64'd354450014208, 64'd33948788736, 64'd2726537728, 64'd73617664, - 64'd371036192768, 64'd32396066816, 64'd2706995200, 64'd75242768, - 64'd386846326784, 64'd30844850176, 64'd2685821696, 64'd76812912, - 64'd401881497600, 64'd29296365568, 64'd2663046912, 64'd78326888, - 64'd416143343616, 64'd27751819264, 64'd2638700544, 64'd79783560, - 64'd429634158592, 64'd26212401152, 64'd2612814336, 64'd81181848, - 64'd442356793344, 64'd24679286784, 64'd2585420544, 64'd82520744, - 64'd454314688512, 64'd23153633280, 64'd2556553472, 64'd83799312, - 64'd465511874560, 64'd21636573184, 64'd2526247424, 64'd85016672, - 64'd475952873472, 64'd20129226752, 64'd2494538240, 64'd86172024, - 64'd485642895360, 64'd18632689664, 64'd2461462784, 64'd87264632, - 64'd494587543552, 64'd17148034048, 64'd2427058944, 64'd88293824, - 64'd502793076736, 64'd15676313600, 64'd2391365376, 64'd89259000, - 64'd510266212352, 64'd14218556416, 64'd2354420992, 64'd90159632, - 64'd517014126592, 64'd12775770112, 64'd2316266496, 64'd90995240, - 64'd523044618240, 64'd11348933632, 64'd2276942592, 64'd91765448, - 64'd528365879296, 64'd9939003392, 64'd2236491264, 64'd92469904, - 64'd532986593280, 64'd8546911744, 64'd2194954752, 64'd93108368, - 64'd536915935232, 64'd7173561856, 64'd2152375552, 64'd93680616, - 64'd540163440640, 64'd5819831808, 64'd2108797824, 64'd94186544, - 64'd542739169280, 64'd4486573056, 64'd2064265216, 64'd94626064, - 64'd544653541376, 64'd3174608640, 64'd2018822272, 64'd94999192, - 64'd545917468672, 64'd1884733568, 64'd1972513664, 64'd95305976, - 64'd546542092288, 64'd617714624, 64'd1925384960, 64'd95546560, - 64'd546539110400, - 64'd625710208, 64'd1877481600, 64'd95721120, - 64'd545920450560, - 64'd1844832128, 64'd1828849408, 64'd95829912, - 64'd544698433536, - 64'd3038971904, 64'd1779534464, 64'd95873240, - 64'd542885740544, - 64'd4207480064, 64'd1729583104, 64'd95851488, - 64'd540495314944, - 64'd5349736960, 64'd1679041664, 64'd95765088, - 64'd537540460544, - 64'd6465153536, 64'd1627956480, 64'd95614512, - 64'd534034743296, - 64'd7553170944, 64'd1576374400, 64'd95400320, - 64'd529991958528, - 64'd8613261312, 64'd1524341760, 64'd95123112, - 64'd525426229248, - 64'd9644926976, 64'd1471905024, 64'd94783544, - 64'd520351842304, - 64'd10647700480, 64'd1419110784, 64'd94382320, - 64'd514783412224, - 64'd11621147648, 64'd1366005120, 64'd93920200, - 64'd508735651840, - 64'd12564862976, 64'd1312634368, 64'd93398000, - 64'd502223568896, - 64'd13478472704, 64'd1259044096, 64'd92816584, - 64'd495262269440, - 64'd14361633792, 64'd1205280256, 64'd92176856, - 64'd487867056128, - 64'd15214034944, 64'd1151388032, 64'd91479784, - 64'd480053395456, - 64'd16035394560, 64'd1097412480, 64'd90726352, - 64'd471836884992, - 64'd16825462784, 64'd1043398272, 64'd89917624, - 64'd463233187840, - 64'd17584019456, 64'd989389632, 64'd89054672, - 64'd454258130944, - 64'd18310875136, 64'd935430336, 64'd88138632, - 64'd444927606784, - 64'd19005870080, 64'd881563648, 64'd87170672, - 64'd435257606144, - 64'd19668875264, 64'd827832448, 64'd86152000, - 64'd425264087040, - 64'd20299794432, 64'd774278848, 64'd85083856, - 64'd414963171328, - 64'd20898553856, 64'd720944576, 64'd83967520, - 64'd404370915328, - 64'd21465116672, 64'd667870656, 64'd82804296, - 64'd393503408128, - 64'd21999468544, 64'd615097408, 64'd81595528, - 64'd382376804352, - 64'd22501629952, 64'd562664512, 64'd80342592, - 64'd371007160320, - 64'd22971641856, 64'd510611008, 64'd79046888, - 64'd359410499584, - 64'd23409582080, 64'd458975104, 64'd77709832, - 64'd347602878464, - 64'd23815548928, 64'd407794272, 64'd76332888, - 64'd335600254976, - 64'd24189671424, 64'd357105184, 64'd74917520, - 64'd323418488832, - 64'd24532105216, 64'd306943680, 64'd73465224, - 64'd311073406976, - 64'd24843030528, 64'd257344752, 64'd71977528, - 64'd298580672512, - 64'd25122652160, 64'd208342576, 64'd70455960, - 64'd285955948544, - 64'd25371203584, 64'd159970368, 64'd68902072, - 64'd273214619648, - 64'd25588940800, 64'd112260464, 64'd67317424, - 64'd260372086784, - 64'd25776146432, 64'd65244268, 64'd65703596, - 64'd247443505152, - 64'd25933123584, 64'd18952236, 64'd64062188, - 64'd234443948032, - 64'd26060197888, - 64'd26586158, 64'd62394792, - 64'd221388242944, - 64'd26157721600, - 64'd71342424, 64'd60703024, - 64'd208291086336, - 64'd26226067456, - 64'd115289064, 64'd58988492, - 64'd195166978048, - 64'd26265624576, - 64'd158399616, 64'd57252828, - 64'd182030188544, - 64'd26276810752, - 64'd200648608, 64'd55497648, - 64'd168894824448, - 64'd26260058112, - 64'd242011664, 64'd53724580, - 64'd155774713856, - 64'd26215821312, - 64'd282465440, 64'd51935256, - 64'd142683504640, - 64'd26144571392, - 64'd321987616, 64'd50131300, - 64'd129634557952, - 64'd26046797824, - 64'd360556992, 64'd48314332, - 64'd116641038336, - 64'd25923008512, - 64'd398153440, 64'd46485976, - 64'd103715799040, - 64'd25773729792, - 64'd434757920, 64'd44647844, - 64'd90871463936, - 64'd25599500288, - 64'd470352448, 64'd42801540, - 64'd78120370176, - 64'd25400875008, - 64'd504920192, 64'd40948668, - 64'd65474560000, - 64'd25178427392, - 64'd538445376, 64'd39090812, - 64'd52945813504, - 64'd24932741120, - 64'd570913344, 64'd37229548, - 64'd40545595392, - 64'd24664412160, - 64'd602310528, 64'd35366440, - 64'd28285073408, - 64'd24374052864, - 64'd632624512, 64'd33503040, - 64'd16175110144, - 64'd24062283776, - 64'd661843904, 64'd31640880, - 64'd4226252032, - 64'd23729739776, - 64'd689958528, 64'd29781480, 64'd7551273984, - 64'd23377063936, - 64'd716959168, 64'd27926338, 64'd19147565056, - 64'd23004909568, - 64'd742837760, 64'd26076936, 64'd30553047040, - 64'd22613938176, - 64'd767587328, 64'd24234734, 64'd41758478336, - 64'd22204823552, - 64'd791202048, 64'd22401170, 64'd52754960384, - 64'd21778241536, - 64'd813677120, 64'd20577660, 64'd63533924352, - 64'd21334876160, - 64'd835008704, 64'd18765600, 64'd74087153664, - 64'd20875419648, - 64'd855194176, 64'd16966354, 64'd84406779904, - 64'd20400570368, - 64'd874231936, 64'd15181266, 64'd94485274624, - 64'd19911026688, - 64'd892121408, 64'd13411651, 64'd104315469824, - 64'd19407495168, - 64'd908862912, 64'd11658797, 64'd113890557952, - 64'd18890684416, - 64'd924457984, 64'd9923964, 64'd123204067328, - 64'd18361305088, - 64'd938909120, 64'd8208380, 64'd132249886720, - 64'd17820069888, - 64'd952219648, 64'd6513247, 64'd141022281728, - 64'd17267693568, - 64'd964394112, 64'd4839731, 64'd149515845632, - 64'd16704888832, - 64'd975437760, 64'd3188970, 64'd157725540352, - 64'd16132372480, - 64'd985357056, 64'd1562069, 64'd165646712832, - 64'd15550857216, - 64'd994159104, - 64'd39902, 64'd173275021312, - 64'd14961054720, - 64'd1001852224, - 64'd1615906, 64'd180606500864, - 64'd14363675648, - 64'd1008445312, - 64'd3164939, 64'd187637547008, - 64'd13759428608, - 64'd1013948352, - 64'd4686034, 64'd194364899328, - 64'd13149016064, - 64'd1018372160, - 64'd6178258, 64'd200785657856, - 64'd12533139456, - 64'd1021728256, - 64'd7640716, 64'd206897250304, - 64'd11912493056, - 64'd1024029120, - 64'd9072546, 64'd212697464832, - 64'd11287769088, - 64'd1025287936, - 64'd10472925, 64'd218184450048, - 64'd10659650560, - 64'd1025518720, - 64'd11841068, 64'd223356665856, - 64'd10028817408, - 64'd1024736192, - 64'd13176226, 64'd228212932608, - 64'd9395940352, - 64'd1022955776, - 64'd14477687, 64'd232752381952, - 64'd8761683968, - 64'd1020193664, - 64'd15744778, 64'd236974489600, - 64'd8126705152, - 64'd1016466752, - 64'd16976866, 64'd240879075328, - 64'd7491652096, - 64'd1011792384, - 64'd18173352, 64'd244466237440, - 64'd6857163264, - 64'd1006188864, - 64'd19333680, 64'd247736434688, - 64'd6223868928, - 64'd999674816, - 64'd20457330, 64'd250690404352, - 64'd5592388608, - 64'd992269568, - 64'd21543820, 64'd253329227776, - 64'd4963332608, - 64'd983993088, - 64'd22592710, 64'd255654248448, - 64'd4337299456, - 64'd974865728, - 64'd23603594, 64'd257667121152, - 64'd3714877184, - 64'd964908416, - 64'd24576108, 64'd259369828352, - 64'd3096642048, - 64'd954142592, - 64'd25509924, 64'd260764565504, - 64'd2483158272, - 64'd942590080, - 64'd26404754, 64'd261853855744, - 64'd1874978048, - 64'd930273216, - 64'd27260348, 64'd262640517120, - 64'd1272640384, - 64'd917214656, - 64'd28076494, 64'd263127564288, - 64'd676671872, - 64'd903437632, - 64'd28853018, 64'd263318339584, - 64'd87585424, - 64'd888965376, - 64'd29589780, 64'd263216381952, 64'd494119680, - 64'd873821888, - 64'd30286680, 64'd262825525248, 64'd1067958016, - 64'd858031040, - 64'd30943656, 64'd262149816320, 64'd1633458304, - 64'd841617344, - 64'd31560682, 64'd261193531392, 64'd2190163968, - 64'd824605312, - 64'd32137764, 64'd259961192448, 64'd2737633280, - 64'd807019840, - 64'd32674948, 64'd258457501696, 64'd3275438592, - 64'd788885952, - 64'd33172316, 64'd256687423488, 64'd3803168512, - 64'd770228800, - 64'd33629976, 64'd254656086016, 64'd4320425984, - 64'd751073856, - 64'd34048084, 64'd252368814080, 64'd4826830848, - 64'd731446464, - 64'd34426820, 64'd249831129088, 64'd5322016768, - 64'd711372288, - 64'd34766396, 64'd247048716288, 64'd5805634560, - 64'd690876992, - 64'd35067064, 64'd244027473920, 64'd6277350912, - 64'd669986240, - 64'd35329100, 64'd240773414912, 64'd6736847872, - 64'd648725760, - 64'd35552820, 64'd237292716032, 64'd7183823872, - 64'd627121344, - 64'd35738560, 64'd233591717888, 64'd7617994240, - 64'd605198656, - 64'd35886692, 64'd229676892160, 64'd8039089664, - 64'd582983360, - 64'd35997620, 64'd225554857984, 64'd8446857728, - 64'd560501120, - 64'd36071772, 64'd221232300032, 64'd8841062400, - 64'd537777344, - 64'd36109608, 64'd216716083200, 64'd9221482496, - 64'd514837408, - 64'd36111604, 64'd212013154304, 64'd9587915776, - 64'd491706656, - 64'd36078280, 64'd207130525696, 64'd9940173824, - 64'd468410144, - 64'd36010168, 64'd202075373568, 64'd10278087680, - 64'd444972768, - 64'd35907824, 64'd196854857728, 64'd10601500672, - 64'd421419264, - 64'd35771840, 64'd191476301824, 64'd10910274560, - 64'd397774112, - 64'd35602824, 64'd185947045888, 64'd11204287488, - 64'd374061536, - 64'd35401396, 64'd180274495488, 64'd11483432960, - 64'd350305568, - 64'd35168220, 64'd174466105344, 64'd11747620864, - 64'd326529888, - 64'd34903956, 64'd168529379328, 64'd11996775424, - 64'd302757952, - 64'd34609308, 64'd162471854080, 64'd12230838272, - 64'd279012800, - 64'd34284976, 64'd156301066240, 64'd12449766400, - 64'd255317248, - 64'd33931692, 64'd150024601600, 64'd12653530112, - 64'd231693680, - 64'd33550202, 64'd143650062336, 64'd12842118144, - 64'd208164128, - 64'd33141266, 64'd137185017856, 64'd13015530496, - 64'd184750272, - 64'd32705664, 64'd130637062144, 64'd13173785600, - 64'd161473392, - 64'd32244184, 64'd124013756416, 64'd13316914176, - 64'd138354304, - 64'd31757632, 64'd117322661888, 64'd13444962304, - 64'd115413440, - 64'd31246826, 64'd110571298816, 64'd13557988352, - 64'd92670792, - 64'd30712592, 64'd103767162880, 64'd13656068096, - 64'd70145880, - 64'd30155772, 64'd96917708800, 64'd13739287552, - 64'd47857776, - 64'd29577214, 64'd90030333952, 64'd13807748096, - 64'd25825048, - 64'd28977778, 64'd83112402944, 64'd13861564416, - 64'd4065793, - 64'd28358328, 64'd76171190272, 64'd13900861440, 64'd17402396, - 64'd27719738, 64'd69213937664, 64'd13925779456, 64'd38562440, - 64'd27062890, 64'd62247784448, 64'd13936468992, 64'd59397776, - 64'd26388666, 64'd55279808512, 64'd13933095936, 64'd79892376, - 64'd25697958, 64'd48317001728, 64'd13915833344, 64'd100030752, - 64'd24991658, 64'd41366261760, 64'd13884868608, 64'd119797944, - 64'd24270660, 64'd34434383872, 64'd13840399360, 64'd139179568, - 64'd23535864, 64'd27528077312, 64'd13782632448, 64'd158161776, - 64'd22788168, 64'd20653932544, 64'd13711788032, 64'd176731296, - 64'd22028472, 64'd13818431488, 64'd13628093440, 64'd194875424, - 64'd21257672, 64'd7027940352, 64'd13531788288, 64'd212582048, - 64'd20476664, 64'd288703872, 64'd13423118336, 64'd229839616, - 64'd19686344, - 64'd6393159680, 64'd13302340608, 64'd246637136, - 64'd18887604, - 64'd13011662848, 64'd13169720320, 64'd262964256, - 64'd18081328, - 64'd19560951808, 64'd13025530880, 64'd278811168, - 64'd17268400, - 64'd26035312640, 64'd12870052864, 64'd294168672, - 64'd16449699, - 64'd32429170688, 64'd12703575040, 64'd309028160, - 64'd15626094, - 64'd38737104896, 64'd12526392320, 64'd323381600, - 64'd14798449, - 64'd44953829376, 64'd12338807808, 64'd337221536, - 64'd13967621, - 64'd51074228224, 64'd12141129728, 64'd350541152, - 64'd13134456, - 64'd57093328896, 64'd11933672448, 64'd363334208, - 64'd12299796, - 64'd63006322688, 64'd11716757504, 64'd375595008, - 64'd11464468, - 64'd68808564736, 64'd11490709504, 64'd387318496, - 64'd10629291, - 64'd74495565824, 64'd11255858176, 64'd398500160, - 64'd9795073, - 64'd80063012864, 64'd11012540416, 64'd409136096, - 64'd8962611, - 64'd85506752512, 64'd10761092096, 64'd419222944, - 64'd8132689, - 64'd90822803456, 64'd10501858304, 64'd428757984, - 64'd7306078, - 64'd96007372800, 64'd10235184128, 64'd437738944, - 64'd6483536};
endpackage
`endif
