`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam N = 1;
	localparam M = 1;
	localparam real Lfr[0:0] = {0.87730575};
	localparam real Lfi[0:0] = {0.0};
	localparam real Lbr[0:0] = {0.87730575};
	localparam real Lbi[0:0] = {0.0};
	localparam real Wfr[0:0] = {-0.1308997};
	localparam real Wfi[0:0] = {-0.0};
	localparam real Wbr[0:0] = {0.1308997};
	localparam real Wbi[0:0] = {0.0};
	localparam real Ffr[0:0][0:19] = '{
		'{-0.46865743, -0.41115588, -0.36070943, -0.31645244, -0.27762556, -0.2435625, -0.21367879, -0.18746164, -0.16446118, -0.14428274, -0.12658007, -0.111049436, -0.09742431, -0.08547091, -0.07498412, -0.065784, -0.057712685, -0.050631672, -0.044419456, -0.038969446}};
	localparam real Ffi[0:0][0:19] = '{
		'{0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0}};
	localparam real Fbr[0:0][0:19] = '{
		'{0.46865743, 0.41115588, 0.36070943, 0.31645244, 0.27762556, 0.2435625, 0.21367879, 0.18746164, 0.16446118, 0.14428274, 0.12658007, 0.111049436, 0.09742431, 0.08547091, 0.07498412, 0.065784, 0.057712685, 0.050631672, 0.044419456, 0.038969446}};
	localparam real Fbi[0:0][0:19] = '{
		'{0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0}};
	localparam real hf[0:299] = {0.061347116, 0.053820178, 0.047216754, 0.04142353, 0.0363411, 0.031882256, 0.02797049, 0.024538672, 0.021527918, 0.018886566, 0.016569294, 0.014536337, 0.012752812, 0.011188116, 0.009815399, 0.008611105, 0.007554573, 0.0066276705, 0.005814493, 0.0051010884, 0.0044752145, 0.0039261314, 0.0034444178, 0.0030218076, 0.0026510493, 0.0023257807, 0.002040421, 0.001790073, 0.0015704414, 0.0013777573, 0.0012087144, 0.0010604121, 0.0009303057, 0.00081616256, 0.00071602414, 0.00062817207, 0.000551099, 0.00048348232, 0.00042416184, 0.00037211963, 0.0003264627, 0.0002864076, 0.00025126705, 0.00022043803, 0.00019339155, 0.00016966353, 0.00014884678, 0.00013058414, 0.00011456222, 0.0001005061, 8.817458e-05, 7.735607e-05, 6.786492e-05, 5.953829e-05, 5.2233285e-05, 4.5824563e-05, 4.0202154e-05, 3.5269582e-05, 3.0942207e-05, 2.7145777e-05, 2.3815146e-05, 2.0893165e-05, 1.8329694e-05, 1.6080747e-05, 1.4107732e-05, 1.2376795e-05, 1.08582335e-05, 9.525991e-06, 8.357207e-06, 7.3318256e-06, 6.432253e-06, 5.6430526e-06, 4.9506825e-06, 4.3432624e-06, 3.8103692e-06, 3.342859e-06, 2.9327093e-06, 2.5728827e-06, 2.2572049e-06, 1.980259e-06, 1.7372926e-06, 1.5241368e-06, 1.337134e-06, 1.1730754e-06, 1.0291458e-06, 9.0287557e-07, 7.920979e-07, 6.949121e-07, 6.096504e-07, 5.348498e-07, 4.6922682e-07, 4.1165538e-07, 3.6114764e-07, 3.1683692e-07, 2.7796284e-07, 2.438584e-07, 2.1393839e-07, 1.8768938e-07, 1.6466099e-07, 1.4445803e-07, 1.2673387e-07, 1.1118435e-07, 9.7542674e-08, 8.557475e-08, 7.507522e-08, 6.586392e-08, 5.77828e-08, 5.0693185e-08, 4.4473424e-08, 3.901679e-08, 3.4229654e-08, 3.0029874e-08, 2.6345381e-08, 2.3112955e-08, 2.027713e-08, 1.7789242e-08, 1.5606606e-08, 1.3691764e-08, 1.2011864e-08, 1.0538078e-08, 9.245117e-09, 8.110794e-09, 7.1156463e-09, 6.2425975e-09, 5.4766667e-09, 4.8047113e-09, 4.215201e-09, 3.6980201e-09, 3.2442944e-09, 2.8462381e-09, 2.4970213e-09, 2.1906512e-09, 1.9218709e-09, 1.6860684e-09, 1.4791975e-09, 1.2977085e-09, 1.1384872e-09, 9.988014e-10, 8.762542e-10, 7.6874285e-10, 6.744226e-10, 5.916748e-10, 5.190797e-10, 4.553916e-10, 3.995177e-10, 3.5049919e-10, 3.0749495e-10, 2.697671e-10, 2.3666824e-10, 2.076304e-10, 1.8215535e-10, 1.5980595e-10, 1.4019867e-10, 1.229971e-10, 1.0790607e-10, 9.4666615e-11, 8.305157e-11, 7.286162e-11, 6.392192e-11, 5.607907e-11, 4.9198493e-11, 4.316212e-11, 3.7866377e-11, 3.322039e-11, 2.914444e-11, 2.5568585e-11, 2.2431468e-11, 1.9679256e-11, 1.7264724e-11, 1.5146443e-11, 1.3288062e-11, 1.1657693e-11, 1.02273615e-11, 8.972523e-12, 7.871647e-12, 6.905841e-12, 6.058534e-12, 5.3151867e-12, 4.6630443e-12, 4.0909155e-12, 3.5889837e-12, 3.148636e-12, 2.7623166e-12, 2.4233963e-12, 2.1260595e-12, 1.8652044e-12, 1.6363546e-12, 1.4355833e-12, 1.2594455e-12, 1.1049188e-12, 9.693517e-13, 8.5041777e-13, 7.4607643e-13, 6.5453713e-13, 5.742292e-13, 5.037746e-13, 4.4196436e-13, 3.8773788e-13, 3.401647e-13, 2.9842844e-13, 2.61813e-13, 2.2969005e-13, 2.015084e-13, 1.7678449e-13, 1.5509405e-13, 1.360649e-13, 1.1937052e-13, 1.0472445e-13, 9.187537e-14, 8.060279e-14, 7.071329e-14, 6.203718e-14, 5.4425573e-14, 4.774787e-14, 4.1889482e-14, 3.6749883e-14, 3.2240886e-14, 2.8285115e-14, 2.4814694e-14, 2.1770075e-14, 1.9099012e-14, 1.6755674e-14, 1.4699849e-14, 1.2896262e-14, 1.1313966e-14, 9.925807e-15, 8.707968e-15, 7.63955e-15, 6.7022215e-15, 5.8798977e-15, 5.1584683e-15, 4.525554e-15, 3.9702946e-15, 3.4831623e-15, 3.0557984e-15, 2.6808697e-15, 2.3519424e-15, 2.0633725e-15, 1.8102087e-15, 1.5881065e-15, 1.393255e-15, 1.2223107e-15, 1.0723402e-15, 9.407703e-16, 8.2534313e-16, 7.240783e-16, 6.352381e-16, 5.57298e-16, 4.8892076e-16, 4.28933e-16, 3.763054e-16, 3.301349e-16, 2.8962926e-16, 2.5409342e-16, 2.2291763e-16, 1.9556691e-16, 1.7157199e-16, 1.5052109e-16, 1.3205302e-16, 1.1585088e-16, 1.0163664e-16, 8.916641e-17, 7.8226206e-17, 6.8628303e-17, 6.020801e-17, 5.2820832e-17, 4.634002e-17, 4.065437e-17, 3.566631e-17, 3.129026e-17, 2.7451127e-17, 2.4083031e-17, 2.1128183e-17, 1.8535877e-17, 1.6261631e-17, 1.4266422e-17, 1.2516015e-17, 1.0980373e-17, 9.6331436e-18, 8.4512125e-18, 7.414298e-18, 6.5046063e-18, 5.7065284e-18, 5.0063705e-18, 4.3921177e-18, 3.8532302e-18, 3.380461e-18, 2.9656979e-18, 2.6018238e-18, 2.2825952e-18, 2.002534e-18, 1.7568344e-18, 1.5412811e-18, 1.3521748e-18, 1.1862707e-18, 1.0407221e-18, 9.130315e-19, 8.0100784e-19, 7.027288e-19, 6.1650805e-19};
	localparam real hb[0:299] = {0.061347116, 0.053820178, 0.047216754, 0.04142353, 0.0363411, 0.031882256, 0.02797049, 0.024538672, 0.021527918, 0.018886566, 0.016569294, 0.014536337, 0.012752812, 0.011188116, 0.009815399, 0.008611105, 0.007554573, 0.0066276705, 0.005814493, 0.0051010884, 0.0044752145, 0.0039261314, 0.0034444178, 0.0030218076, 0.0026510493, 0.0023257807, 0.002040421, 0.001790073, 0.0015704414, 0.0013777573, 0.0012087144, 0.0010604121, 0.0009303057, 0.00081616256, 0.00071602414, 0.00062817207, 0.000551099, 0.00048348232, 0.00042416184, 0.00037211963, 0.0003264627, 0.0002864076, 0.00025126705, 0.00022043803, 0.00019339155, 0.00016966353, 0.00014884678, 0.00013058414, 0.00011456222, 0.0001005061, 8.817458e-05, 7.735607e-05, 6.786492e-05, 5.953829e-05, 5.2233285e-05, 4.5824563e-05, 4.0202154e-05, 3.5269582e-05, 3.0942207e-05, 2.7145777e-05, 2.3815146e-05, 2.0893165e-05, 1.8329694e-05, 1.6080747e-05, 1.4107732e-05, 1.2376795e-05, 1.08582335e-05, 9.525991e-06, 8.357207e-06, 7.3318256e-06, 6.432253e-06, 5.6430526e-06, 4.9506825e-06, 4.3432624e-06, 3.8103692e-06, 3.342859e-06, 2.9327093e-06, 2.5728827e-06, 2.2572049e-06, 1.980259e-06, 1.7372926e-06, 1.5241368e-06, 1.337134e-06, 1.1730754e-06, 1.0291458e-06, 9.0287557e-07, 7.920979e-07, 6.949121e-07, 6.096504e-07, 5.348498e-07, 4.6922682e-07, 4.1165538e-07, 3.6114764e-07, 3.1683692e-07, 2.7796284e-07, 2.438584e-07, 2.1393839e-07, 1.8768938e-07, 1.6466099e-07, 1.4445803e-07, 1.2673387e-07, 1.1118435e-07, 9.7542674e-08, 8.557475e-08, 7.507522e-08, 6.586392e-08, 5.77828e-08, 5.0693185e-08, 4.4473424e-08, 3.901679e-08, 3.4229654e-08, 3.0029874e-08, 2.6345381e-08, 2.3112955e-08, 2.027713e-08, 1.7789242e-08, 1.5606606e-08, 1.3691764e-08, 1.2011864e-08, 1.0538078e-08, 9.245117e-09, 8.110794e-09, 7.1156463e-09, 6.2425975e-09, 5.4766667e-09, 4.8047113e-09, 4.215201e-09, 3.6980201e-09, 3.2442944e-09, 2.8462381e-09, 2.4970213e-09, 2.1906512e-09, 1.9218709e-09, 1.6860684e-09, 1.4791975e-09, 1.2977085e-09, 1.1384872e-09, 9.988014e-10, 8.762542e-10, 7.6874285e-10, 6.744226e-10, 5.916748e-10, 5.190797e-10, 4.553916e-10, 3.995177e-10, 3.5049919e-10, 3.0749495e-10, 2.697671e-10, 2.3666824e-10, 2.076304e-10, 1.8215535e-10, 1.5980595e-10, 1.4019867e-10, 1.229971e-10, 1.0790607e-10, 9.4666615e-11, 8.305157e-11, 7.286162e-11, 6.392192e-11, 5.607907e-11, 4.9198493e-11, 4.316212e-11, 3.7866377e-11, 3.322039e-11, 2.914444e-11, 2.5568585e-11, 2.2431468e-11, 1.9679256e-11, 1.7264724e-11, 1.5146443e-11, 1.3288062e-11, 1.1657693e-11, 1.02273615e-11, 8.972523e-12, 7.871647e-12, 6.905841e-12, 6.058534e-12, 5.3151867e-12, 4.6630443e-12, 4.0909155e-12, 3.5889837e-12, 3.148636e-12, 2.7623166e-12, 2.4233963e-12, 2.1260595e-12, 1.8652044e-12, 1.6363546e-12, 1.4355833e-12, 1.2594455e-12, 1.1049188e-12, 9.693517e-13, 8.5041777e-13, 7.4607643e-13, 6.5453713e-13, 5.742292e-13, 5.037746e-13, 4.4196436e-13, 3.8773788e-13, 3.401647e-13, 2.9842844e-13, 2.61813e-13, 2.2969005e-13, 2.015084e-13, 1.7678449e-13, 1.5509405e-13, 1.360649e-13, 1.1937052e-13, 1.0472445e-13, 9.187537e-14, 8.060279e-14, 7.071329e-14, 6.203718e-14, 5.4425573e-14, 4.774787e-14, 4.1889482e-14, 3.6749883e-14, 3.2240886e-14, 2.8285115e-14, 2.4814694e-14, 2.1770075e-14, 1.9099012e-14, 1.6755674e-14, 1.4699849e-14, 1.2896262e-14, 1.1313966e-14, 9.925807e-15, 8.707968e-15, 7.63955e-15, 6.7022215e-15, 5.8798977e-15, 5.1584683e-15, 4.525554e-15, 3.9702946e-15, 3.4831623e-15, 3.0557984e-15, 2.6808697e-15, 2.3519424e-15, 2.0633725e-15, 1.8102087e-15, 1.5881065e-15, 1.393255e-15, 1.2223107e-15, 1.0723402e-15, 9.407703e-16, 8.2534313e-16, 7.240783e-16, 6.352381e-16, 5.57298e-16, 4.8892076e-16, 4.28933e-16, 3.763054e-16, 3.301349e-16, 2.8962926e-16, 2.5409342e-16, 2.2291763e-16, 1.9556691e-16, 1.7157199e-16, 1.5052109e-16, 1.3205302e-16, 1.1585088e-16, 1.0163664e-16, 8.916641e-17, 7.8226206e-17, 6.8628303e-17, 6.020801e-17, 5.2820832e-17, 4.634002e-17, 4.065437e-17, 3.566631e-17, 3.129026e-17, 2.7451127e-17, 2.4083031e-17, 2.1128183e-17, 1.8535877e-17, 1.6261631e-17, 1.4266422e-17, 1.2516015e-17, 1.0980373e-17, 9.6331436e-18, 8.4512125e-18, 7.414298e-18, 6.5046063e-18, 5.7065284e-18, 5.0063705e-18, 4.3921177e-18, 3.8532302e-18, 3.380461e-18, 2.9656979e-18, 2.6018238e-18, 2.2825952e-18, 2.002534e-18, 1.7568344e-18, 1.5412811e-18, 1.3521748e-18, 1.1862707e-18, 1.0407221e-18, 9.130315e-19, 8.0100784e-19, 7.027288e-19, 6.1650805e-19};
endpackage
`endif
