`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam N = 4;
	localparam COEFF_BIAS = 48;
	localparam logic signed[63:0] Lfr[0:3] = {64'(277489893271481), 64'(277489893271481), 64'(275315491622285), 64'(275315491622285)};
	localparam logic signed[63:0] Lfi[0:3] = {64'(30020001337947), 64'(-30020001337947), 64'(11558098293529), 64'(-11558098293529)};
	localparam logic signed[63:0] Lbr[0:3] = {64'(277489893271481), 64'(277489893271481), 64'(275315491622285), 64'(275315491622285)};
	localparam logic signed[63:0] Lbi[0:3] = {64'(30020001337947), 64'(-30020001337947), 64'(11558098293529), 64'(-11558098293529)};
	localparam logic signed[63:0] Wfr[0:3] = {64'(24193209882), 64'(24193209882), 64'(-7887428590), 64'(-7887428590)};
	localparam logic signed[63:0] Wfi[0:3] = {64'(29297075841), 64'(-29297075841), 64'(-33126712469), 64'(33126712469)};
	localparam logic signed[63:0] Wbr[0:3] = {64'(-24193209882), 64'(-24193209882), 64'(7887428590), 64'(7887428590)};
	localparam logic signed[63:0] Wbi[0:3] = {64'(-29297075841), 64'(29297075841), 64'(33126712469), 64'(-33126712469)};
	localparam logic signed[63:0] Ffr[0:3][0:79] = '{
		'{64'(2678910912348682), 64'(1633669149297615), 64'(-134405106412023), 64'(-14489081406757), 64'(3471761733289509), 64'(1534935316807140), 64'(-154547576200402), 64'(-12167341321049), 64'(4211153497515380), 64'(1420087166233641), 64'(-172563932222687), 64'(-9743629047954), 64'(4889422534499934), 64'(1290723849399400), 64'(-188281223922595), 64'(-7247706595933), 64'(5499740975037776), 64'(1148585763351890), 64'(-201556008143343), 64'(-4709673588602), 64'(6036181793402482), 64'(995532040410431), 64'(-212275515540637), 64'(-2159613203878), 64'(6493772333226378), 64'(833517040657504), 64'(-220358442413966), 64'(372755769329), 64'(6868535890318197), 64'(664566135678268), 64'(-225755365061278), 64'(2858416831816), 64'(7157521071022570), 64'(490751075721102), 64'(-228448778179966), 64'(5269379888993), 64'(7358818790936519), 64'(314165232382821), 64'(-228452763163329), 64'(7578988059119), 64'(7471566924126414), 64'(136899005473061), 64'(-225812296327788), 64'(9762203913194), 64'(7495942755766966), 64'(-38984324020268), 64'(-220602211106000), 64'(11795872177577), 64'(7433143529741519), 64'(-211472022825834), 64'(-212925832011491), 64'(13658956252499), 64'(7285355515665612), 64'(-378624356972050), 64'(-202913301681643), 64'(15332746247078), 64'(7055712145579892), 64'(-538595822537850), 64'(-190719625501872), 64'(16801036599608), 64'(6748241887867779), 64'(-689654930258371), 64'(-176522461172683), 64'(18050271736293), 64'(6367806633571694), 64'(-830202339184127), 64'(-160519683075600), 64'(19069658617453), 64'(5920031467125635), 64'(-958787157130758), 64'(-142926753400873), 64'(19851245422781), 64'(5411226778650929), 64'(-1074121249927379), 64'(-123973933701595), 64'(20389966031699), 64'(4848303747586724), 64'(-1175091427164946), 64'(-103903371822373), 64'(20683650356549)},
		'{64'(2678910912348222), 64'(1633669149297648), 64'(-134405106412032), 64'(-14489081406755), 64'(3471761733289070), 64'(1534935316807172), 64'(-154547576200411), 64'(-12167341321048), 64'(4211153497514966), 64'(1420087166233671), 64'(-172563932222695), 64'(-9743629047952), 64'(4889422534499551), 64'(1290723849399429), 64'(-188281223922603), 64'(-7247706595932), 64'(5499740975037427), 64'(1148585763351916), 64'(-201556008143349), 64'(-4709673588600), 64'(6036181793402171), 64'(995532040410455), 64'(-212275515540643), 64'(-2159613203877), 64'(6493772333226108), 64'(833517040657526), 64'(-220358442413972), 64'(372755769330), 64'(6868535890317968), 64'(664566135678286), 64'(-225755365061283), 64'(2858416831817), 64'(7157521071022387), 64'(490751075721118), 64'(-228448778179969), 64'(5269379888994), 64'(7358818790936382), 64'(314165232382833), 64'(-228452763163332), 64'(7578988059119), 64'(7471566924126326), 64'(136899005473070), 64'(-225812296327790), 64'(9762203913194), 64'(7495942755766923), 64'(-38984324020262), 64'(-220602211106001), 64'(11795872177577), 64'(7433143529741523), 64'(-211472022825831), 64'(-212925832011491), 64'(13658956252499), 64'(7285355515665663), 64'(-378624356972050), 64'(-202913301681642), 64'(15332746247078), 64'(7055712145579987), 64'(-538595822537854), 64'(-190719625501870), 64'(16801036599608), 64'(6748241887867917), 64'(-689654930258378), 64'(-176522461172680), 64'(18050271736292), 64'(6367806633571872), 64'(-830202339184137), 64'(-160519683075597), 64'(19069658617452), 64'(5920031467125852), 64'(-958787157130771), 64'(-142926753400869), 64'(19851245422781), 64'(5411226778651180), 64'(-1074121249927394), 64'(-123973933701590), 64'(20389966031698), 64'(4848303747587006), 64'(-1175091427164964), 64'(-103903371822367), 64'(20683650356548)},
		'{64'(-2621464726625032), 64'(-1601298142322358), 64'(114277463862052), 64'(-54557765512014), 64'(-3402192470904109), 64'(-1521613693668172), 64'(101035526953527), 64'(-52555428834631), 64'(-4143075592769200), 64'(-1441949887694716), 64'(88125723066021), 64'(-50522608463608), 64'(-4844167648167600), 64'(-1362478337710847), 64'(75562184921028), 64'(-48464973598293), 64'(-5505606112696863), 64'(-1283363101544773), 64'(63357707642890), 64'(-46388011318305), 64'(-6127608592847788), 64'(-1204760640672868), 64'(51523776702445), 64'(-44297022280332), 64'(-6710469021379336), 64'(-1126819797494854), 64'(40070597533593), 64'(-42197116997554), 64'(-7254553845722606), 64'(-1049681790049648), 64'(29007126689070), 64'(-40093212685504), 64'(-7760298217955961), 64'(-973480223457764), 64'(18341104403946), 64'(-37990030657633), 64'(-8228202194534652), 64'(-898341117369665), 64'(8079088437780), 64'(-35892094253348), 64'(-8658826953596720), 64'(-824382948694780), 64'(-1773510931025), 64'(-33803727280864), 64'(-9052791037303526), 64'(-751716708882984), 64'(-11212394882364), 64'(-31729052956814), 64'(-9410766626308762), 64'(-680445975029133), 64'(-20234339123843), 64'(-29671993324251), 64'(-9733475853085184), 64'(-610666994071677), 64'(-28837156170190), 64'(-27636269130411), 64'(-10021687160474126), 64'(-542468779358319), 64'(-37019656947170), 64'(-25625400145358), 64'(-10276211711460314), 64'(-475933218855185), 64'(-44781611831263), 64'(-23642705902492), 64'(-10497899855813746), 64'(-411135194280852), 64'(-52123711232903), 64'(-21691306841762), 64'(-10687637658882664), 64'(-348142710452834), 64'(-59047525827614), 64'(-19774125836360), 64'(-10846343497467206), 64'(-287017034141629), 64'(-65555466535792), 64'(-17893890083631), 64'(-10974964727353150), 64'(-227812841736200), 64'(-71650744348225), 64'(-16053133340965)},
		'{64'(-2621464726623828), 64'(-1601298142322414), 64'(114277463862073), 64'(-54557765512018), 64'(-3402192470902937), 64'(-1521613693668227), 64'(101035526953548), 64'(-52555428834635), 64'(-4143075592768060), 64'(-1441949887694769), 64'(88125723066041), 64'(-50522608463611), 64'(-4844167648166494), 64'(-1362478337710898), 64'(75562184921047), 64'(-48464973598296), 64'(-5505606112695792), 64'(-1283363101544822), 64'(63357707642909), 64'(-46388011318308), 64'(-6127608592846752), 64'(-1204760640672916), 64'(51523776702463), 64'(-44297022280336), 64'(-6710469021378337), 64'(-1126819797494900), 64'(40070597533610), 64'(-42197116997558), 64'(-7254553845721645), 64'(-1049681790049693), 64'(29007126689086), 64'(-40093212685508), 64'(-7760298217955038), 64'(-973480223457806), 64'(18341104403961), 64'(-37990030657636), 64'(-8228202194533767), 64'(-898341117369706), 64'(8079088437795), 64'(-35892094253351), 64'(-8658826953595873), 64'(-824382948694820), 64'(-1773510931011), 64'(-33803727280867), 64'(-9052791037302716), 64'(-751716708883021), 64'(-11212394882350), 64'(-31729052956816), 64'(-9410766626307994), 64'(-680445975029168), 64'(-20234339123830), 64'(-29671993324253), 64'(-9733475853084454), 64'(-610666994071711), 64'(-28837156170178), 64'(-27636269130413), 64'(-10021687160473434), 64'(-542468779358351), 64'(-37019656947158), 64'(-25625400145361), 64'(-10276211711459662), 64'(-475933218855215), 64'(-44781611831252), 64'(-23642705902494), 64'(-10497899855813134), 64'(-411135194280880), 64'(-52123711232892), 64'(-21691306841764), 64'(-10687637658882086), 64'(-348142710452861), 64'(-59047525827604), 64'(-19774125836362), 64'(-10846343497466668), 64'(-287017034141654), 64'(-65555466535783), 64'(-17893890083633), 64'(-10974964727352650), 64'(-227812841736223), 64'(-71650744348217), 64'(-16053133340967)}};
	localparam logic signed[63:0] Ffi[0:3][0:79] = '{
		'{64'(-7789584925020542), 64'(708887221199158), 64'(206702748225345), 64'(-19845819841343), 64'(-7393588604643268), 64'(873085743790186), 64'(189441643064671), 64'(-21110141804839), 64'(-6918639246994867), 64'(1024429359565470), 64'(170276674079435), 64'(-22108944360993), 64'(-6371556198568730), 64'(1161381434685642), 64'(149461551191332), 64'(-22835111110926), 64'(-5759879607888508), 64'(1282597644249564), 64'(127264837936302), 64'(-23284800600437), 64'(-5091771080218742), 64'(1386938313763277), 64'(103966594132111), 64'(-23457435961284), 64'(-4375908801885497), 64'(1473478185138040), 64'(79854941677750), 64'(-23355656937657), 64'(-3621378440744956), 64'(1541513537288885), 64'(55222594523002), 64'(-22985235482842), 64'(-2837561156357778), 64'(1590566623196748), 64'(30363393574268), 64'(-22354956512906), 64'(-2034020064558232), 64'(1620387416998140), 64'(5568886563156), 64'(-21476465781011), 64'(-1220386496487038), 64'(1630952695911008), 64'(-18875008286193), 64'(-20364087183631), 64'(-406247372102465), 64'(1622462512239921), 64'(-42691217575166), 64'(-19034612125145), 64'(398965026813756), 64'(1595334139989243), 64'(-65614571842042), 64'(-17507063846684), 64'(1186079648425665), 64'(1550193608429831), 64'(-87394675671855), 64'(-15802439866300), 64'(1946288454422587), 64'(1487864961015521), 64'(-107798558746626), 64'(-13943435878179), 64'(2671242297735851), 64'(1409357402058381), 64'(-126613080816752), 64'(-11954154617209), 64'(3353139883456778), 64'(1315850515302490), 64'(-143647066875003), 64'(-9859803310541), 64'(3984808899006887), 64'(1208677757771555), 64'(-158733152334642), 64'(-7686383409257), 64'(4559778505553668), 64'(1089308448825112), 64'(-171729321708043), 64'(-5460376320793), 64'(5072342496187033), 64'(959328488094488), 64'(-182520128106280), 64'(-3208428846785)},
		'{64'(7789584925020678), 64'(-708887221199165), 64'(-206702748225342), 64'(19845819841342), 64'(7393588604643451), 64'(-873085743790196), 64'(-189441643064668), 64'(21110141804838), 64'(6918639246995094), 64'(-1024429359565484), 64'(-170276674079431), 64'(22108944360992), 64'(6371556198568998), 64'(-1161381434685658), 64'(-149461551191327), 64'(22835111110925), 64'(5759879607888814), 64'(-1282597644249583), 64'(-127264837936296), 64'(23284800600436), 64'(5091771080219080), 64'(-1386938313763298), 64'(-103966594132105), 64'(23457435961283), 64'(4375908801885863), 64'(-1473478185138064), 64'(-79854941677743), 64'(23355656937656), 64'(3621378440745346), 64'(-1541513537288910), 64'(-55222594522994), 64'(22985235482840), 64'(2837561156358186), 64'(-1590566623196775), 64'(-30363393574260), 64'(22354956512905), 64'(2034020064558654), 64'(-1620387416998168), 64'(-5568886563148), 64'(21476465781009), 64'(1220386496487468), 64'(-1630952695911038), 64'(18875008286202), 64'(20364087183629), 64'(406247372102900), 64'(-1622462512239951), 64'(42691217575174), 64'(19034612125143), 64'(-398965026813322), 64'(-1595334139989273), 64'(65614571842050), 64'(17507063846682), 64'(-1186079648425238), 64'(-1550193608429861), 64'(87394675671863), 64'(15802439866299), 64'(-1946288454422172), 64'(-1487864961015550), 64'(107798558746634), 64'(13943435878177), 64'(-2671242297735452), 64'(-1409357402058410), 64'(126613080816760), 64'(11954154617207), 64'(-3353139883456400), 64'(-1315850515302518), 64'(143647066875011), 64'(9859803310540), 64'(-3984808899006532), 64'(-1208677757771581), 64'(158733152334649), 64'(7686383409256), 64'(-4559778505553342), 64'(-1089308448825137), 64'(171729321708049), 64'(5460376320792), 64'(-5072342496186738), 64'(-959328488094511), 64'(182520128106285), 64'(3208428846784)},
		'{64'(20410122023596984), 64'(-1087203619517777), 64'(261581401330405), 64'(-19688353631198), 64'(19855845437227768), 64'(-1129165953014674), 64'(260549776479662), 64'(-21497800075813), 64'(19281639300793944), 64'(-1166937977762846), 64'(258996978016206), 64'(-23185429430581), 64'(18689575854732616), 64'(-1200612237457261), 64'(256948048973282), 64'(-24752655664962), 64'(18081679793730520), 64'(-1230286297560720), 64'(254428064696757), 64'(-26201094598827), 64'(17459925861202104), 64'(-1256062325165291), 64'(251462077212791), 64'(-27532552007075), 64'(16826236651983674), 64'(-1278046676369314), 64'(248075061960339), 64'(-28749011807856), 64'(16182480619338714), 64'(-1296349491750649), 64'(244291866905447), 64'(-29852624356494), 64'(15530470282089826), 64'(-1311084300475151), 64'(240137164048391), 64'(-30845694866052), 64'(14871960627433400), 64'(-1322367633538259), 64'(235635403329143), 64'(-31730671974348), 64'(14208647704754270), 64'(-1330318646597064), 64'(230810768931151), 64'(-32510136476076), 64'(13542167405539158), 64'(-1335058752810478), 64'(225687137978284), 64'(-33186790237559), 64'(12874094424288384), 64'(-1336711266066034), 64'(220288041614798), 64'(-33763445310536), 64'(12205941395145922), 64'(-1335401054933668), 64'(214636628453457), 64'(-34243013260277), 64'(11539158198806890), 64'(-1331254207649389), 64'(208755630372409), 64'(-34628494722203), 64'(10875131434119388), 64'(-1324397708395326), 64'(202667330637182), 64'(-34922969200132), 64'(10215184048673250), 64'(-1314959125107046), 64'(196393534320064), 64'(-35129585118164), 64'(9560575122561506), 64'(-1303066309004502), 64'(189955540985356), 64'(-35251550137213), 64'(8912499799410572), 64'(-1288847106009427), 64'(183374119605357), 64'(-35292121746123), 64'(8272089358702066), 64'(-1272429080179444), 64'(176669485668604), 64'(-35254598136332)},
		'{64'(-20410122023597112), 64'(1087203619517783), 64'(-261581401330408), 64'(19688353631199), 64'(-19855845437227944), 64'(1129165953014683), 64'(-260549776479665), 64'(21497800075814), 64'(-19281639300794168), 64'(1166937977762856), 64'(-258996978016210), 64'(23185429430582), 64'(-18689575854732880), 64'(1200612237457274), 64'(-256948048973287), 64'(24752655664963), 64'(-18081679793730820), 64'(1230286297560734), 64'(-254428064696763), 64'(26201094598828), 64'(-17459925861202444), 64'(1256062325165307), 64'(-251462077212797), 64'(27532552007076), 64'(-16826236651984046), 64'(1278046676369332), 64'(-248075061960346), 64'(28749011807857), 64'(-16182480619339120), 64'(1296349491750668), 64'(-244291866905454), 64'(29852624356495), 64'(-15530470282090264), 64'(1311084300475172), 64'(-240137164048399), 64'(30845694866053), 64'(-14871960627433864), 64'(1322367633538281), 64'(-235635403329152), 64'(31730671974350), 64'(-14208647704754760), 64'(1330318646597088), 64'(-230810768931160), 64'(32510136476078), 64'(-13542167405539672), 64'(1335058752810502), 64'(-225687137978293), 64'(33186790237561), 64'(-12874094424288920), 64'(1336711266066060), 64'(-220288041614808), 64'(33763445310538), 64'(-12205941395146478), 64'(1335401054933694), 64'(-214636628453467), 64'(34243013260279), 64'(-11539158198807466), 64'(1331254207649416), 64'(-208755630372419), 64'(34628494722205), 64'(-10875131434119980), 64'(1324397708395354), 64'(-202667330637193), 64'(34922969200134), 64'(-10215184048673856), 64'(1314959125107074), 64'(-196393534320075), 64'(35129585118166), 64'(-9560575122562122), 64'(1303066309004531), 64'(-189955540985367), 64'(35251550137215), 64'(-8912499799411199), 64'(1288847106009456), 64'(-183374119605368), 64'(35292121746125), 64'(-8272089358702702), 64'(1272429080179473), 64'(-176669485668615), 64'(35254598136334)}};
	localparam logic signed[63:0] Fbr[0:3][0:79] = '{
		'{64'(-2678910912348682), 64'(1633669149297615), 64'(134405106412023), 64'(-14489081406757), 64'(-3471761733289509), 64'(1534935316807140), 64'(154547576200402), 64'(-12167341321049), 64'(-4211153497515380), 64'(1420087166233641), 64'(172563932222687), 64'(-9743629047954), 64'(-4889422534499934), 64'(1290723849399400), 64'(188281223922595), 64'(-7247706595933), 64'(-5499740975037776), 64'(1148585763351890), 64'(201556008143343), 64'(-4709673588602), 64'(-6036181793402482), 64'(995532040410431), 64'(212275515540637), 64'(-2159613203878), 64'(-6493772333226378), 64'(833517040657504), 64'(220358442413966), 64'(372755769329), 64'(-6868535890318197), 64'(664566135678268), 64'(225755365061278), 64'(2858416831816), 64'(-7157521071022570), 64'(490751075721102), 64'(228448778179966), 64'(5269379888993), 64'(-7358818790936519), 64'(314165232382821), 64'(228452763163329), 64'(7578988059119), 64'(-7471566924126414), 64'(136899005473061), 64'(225812296327788), 64'(9762203913194), 64'(-7495942755766966), 64'(-38984324020268), 64'(220602211106000), 64'(11795872177577), 64'(-7433143529741519), 64'(-211472022825834), 64'(212925832011491), 64'(13658956252499), 64'(-7285355515665612), 64'(-378624356972050), 64'(202913301681643), 64'(15332746247078), 64'(-7055712145579892), 64'(-538595822537850), 64'(190719625501872), 64'(16801036599608), 64'(-6748241887867779), 64'(-689654930258371), 64'(176522461172683), 64'(18050271736293), 64'(-6367806633571694), 64'(-830202339184127), 64'(160519683075600), 64'(19069658617453), 64'(-5920031467125635), 64'(-958787157130758), 64'(142926753400873), 64'(19851245422781), 64'(-5411226778650929), 64'(-1074121249927379), 64'(123973933701595), 64'(20389966031699), 64'(-4848303747586724), 64'(-1175091427164946), 64'(103903371822373), 64'(20683650356549)},
		'{64'(-2678910912348222), 64'(1633669149297648), 64'(134405106412032), 64'(-14489081406755), 64'(-3471761733289070), 64'(1534935316807172), 64'(154547576200411), 64'(-12167341321048), 64'(-4211153497514966), 64'(1420087166233671), 64'(172563932222695), 64'(-9743629047952), 64'(-4889422534499551), 64'(1290723849399429), 64'(188281223922603), 64'(-7247706595932), 64'(-5499740975037427), 64'(1148585763351916), 64'(201556008143349), 64'(-4709673588600), 64'(-6036181793402171), 64'(995532040410455), 64'(212275515540643), 64'(-2159613203877), 64'(-6493772333226108), 64'(833517040657526), 64'(220358442413972), 64'(372755769330), 64'(-6868535890317968), 64'(664566135678286), 64'(225755365061283), 64'(2858416831817), 64'(-7157521071022387), 64'(490751075721118), 64'(228448778179969), 64'(5269379888994), 64'(-7358818790936382), 64'(314165232382833), 64'(228452763163332), 64'(7578988059119), 64'(-7471566924126326), 64'(136899005473070), 64'(225812296327790), 64'(9762203913194), 64'(-7495942755766923), 64'(-38984324020262), 64'(220602211106001), 64'(11795872177577), 64'(-7433143529741523), 64'(-211472022825831), 64'(212925832011491), 64'(13658956252499), 64'(-7285355515665663), 64'(-378624356972050), 64'(202913301681642), 64'(15332746247078), 64'(-7055712145579987), 64'(-538595822537854), 64'(190719625501870), 64'(16801036599608), 64'(-6748241887867917), 64'(-689654930258378), 64'(176522461172680), 64'(18050271736292), 64'(-6367806633571872), 64'(-830202339184137), 64'(160519683075597), 64'(19069658617452), 64'(-5920031467125852), 64'(-958787157130771), 64'(142926753400869), 64'(19851245422781), 64'(-5411226778651180), 64'(-1074121249927394), 64'(123973933701590), 64'(20389966031698), 64'(-4848303747587006), 64'(-1175091427164964), 64'(103903371822367), 64'(20683650356548)},
		'{64'(2621464726625032), 64'(-1601298142322358), 64'(-114277463862052), 64'(-54557765512014), 64'(3402192470904109), 64'(-1521613693668172), 64'(-101035526953527), 64'(-52555428834631), 64'(4143075592769200), 64'(-1441949887694716), 64'(-88125723066021), 64'(-50522608463608), 64'(4844167648167600), 64'(-1362478337710847), 64'(-75562184921028), 64'(-48464973598293), 64'(5505606112696863), 64'(-1283363101544773), 64'(-63357707642890), 64'(-46388011318305), 64'(6127608592847788), 64'(-1204760640672868), 64'(-51523776702445), 64'(-44297022280332), 64'(6710469021379336), 64'(-1126819797494854), 64'(-40070597533593), 64'(-42197116997554), 64'(7254553845722606), 64'(-1049681790049648), 64'(-29007126689070), 64'(-40093212685504), 64'(7760298217955961), 64'(-973480223457764), 64'(-18341104403946), 64'(-37990030657633), 64'(8228202194534652), 64'(-898341117369665), 64'(-8079088437780), 64'(-35892094253348), 64'(8658826953596720), 64'(-824382948694780), 64'(1773510931025), 64'(-33803727280864), 64'(9052791037303526), 64'(-751716708882984), 64'(11212394882364), 64'(-31729052956814), 64'(9410766626308762), 64'(-680445975029133), 64'(20234339123843), 64'(-29671993324251), 64'(9733475853085184), 64'(-610666994071677), 64'(28837156170190), 64'(-27636269130411), 64'(10021687160474126), 64'(-542468779358319), 64'(37019656947170), 64'(-25625400145358), 64'(10276211711460314), 64'(-475933218855185), 64'(44781611831263), 64'(-23642705902492), 64'(10497899855813746), 64'(-411135194280852), 64'(52123711232903), 64'(-21691306841762), 64'(10687637658882664), 64'(-348142710452834), 64'(59047525827614), 64'(-19774125836360), 64'(10846343497467206), 64'(-287017034141629), 64'(65555466535792), 64'(-17893890083631), 64'(10974964727353150), 64'(-227812841736200), 64'(71650744348225), 64'(-16053133340965)},
		'{64'(2621464726623828), 64'(-1601298142322414), 64'(-114277463862073), 64'(-54557765512018), 64'(3402192470902937), 64'(-1521613693668227), 64'(-101035526953548), 64'(-52555428834635), 64'(4143075592768060), 64'(-1441949887694769), 64'(-88125723066041), 64'(-50522608463611), 64'(4844167648166494), 64'(-1362478337710898), 64'(-75562184921047), 64'(-48464973598296), 64'(5505606112695792), 64'(-1283363101544822), 64'(-63357707642909), 64'(-46388011318308), 64'(6127608592846752), 64'(-1204760640672916), 64'(-51523776702463), 64'(-44297022280336), 64'(6710469021378337), 64'(-1126819797494900), 64'(-40070597533610), 64'(-42197116997558), 64'(7254553845721645), 64'(-1049681790049693), 64'(-29007126689086), 64'(-40093212685508), 64'(7760298217955038), 64'(-973480223457806), 64'(-18341104403961), 64'(-37990030657636), 64'(8228202194533767), 64'(-898341117369706), 64'(-8079088437795), 64'(-35892094253351), 64'(8658826953595873), 64'(-824382948694820), 64'(1773510931011), 64'(-33803727280867), 64'(9052791037302716), 64'(-751716708883021), 64'(11212394882350), 64'(-31729052956816), 64'(9410766626307994), 64'(-680445975029168), 64'(20234339123830), 64'(-29671993324253), 64'(9733475853084454), 64'(-610666994071711), 64'(28837156170178), 64'(-27636269130413), 64'(10021687160473434), 64'(-542468779358351), 64'(37019656947158), 64'(-25625400145361), 64'(10276211711459662), 64'(-475933218855215), 64'(44781611831252), 64'(-23642705902494), 64'(10497899855813134), 64'(-411135194280880), 64'(52123711232892), 64'(-21691306841764), 64'(10687637658882086), 64'(-348142710452861), 64'(59047525827604), 64'(-19774125836362), 64'(10846343497466668), 64'(-287017034141654), 64'(65555466535783), 64'(-17893890083633), 64'(10974964727352650), 64'(-227812841736223), 64'(71650744348217), 64'(-16053133340967)}};
	localparam logic signed[63:0] Fbi[0:3][0:79] = '{
		'{64'(7789584925020542), 64'(708887221199158), 64'(-206702748225345), 64'(-19845819841343), 64'(7393588604643268), 64'(873085743790186), 64'(-189441643064671), 64'(-21110141804839), 64'(6918639246994867), 64'(1024429359565470), 64'(-170276674079435), 64'(-22108944360993), 64'(6371556198568730), 64'(1161381434685642), 64'(-149461551191332), 64'(-22835111110926), 64'(5759879607888508), 64'(1282597644249564), 64'(-127264837936302), 64'(-23284800600437), 64'(5091771080218742), 64'(1386938313763277), 64'(-103966594132111), 64'(-23457435961284), 64'(4375908801885497), 64'(1473478185138040), 64'(-79854941677750), 64'(-23355656937657), 64'(3621378440744956), 64'(1541513537288885), 64'(-55222594523002), 64'(-22985235482842), 64'(2837561156357778), 64'(1590566623196748), 64'(-30363393574268), 64'(-22354956512906), 64'(2034020064558232), 64'(1620387416998140), 64'(-5568886563156), 64'(-21476465781011), 64'(1220386496487038), 64'(1630952695911008), 64'(18875008286193), 64'(-20364087183631), 64'(406247372102465), 64'(1622462512239921), 64'(42691217575166), 64'(-19034612125145), 64'(-398965026813756), 64'(1595334139989243), 64'(65614571842042), 64'(-17507063846684), 64'(-1186079648425665), 64'(1550193608429831), 64'(87394675671855), 64'(-15802439866300), 64'(-1946288454422587), 64'(1487864961015521), 64'(107798558746626), 64'(-13943435878179), 64'(-2671242297735851), 64'(1409357402058381), 64'(126613080816752), 64'(-11954154617209), 64'(-3353139883456778), 64'(1315850515302490), 64'(143647066875003), 64'(-9859803310541), 64'(-3984808899006887), 64'(1208677757771555), 64'(158733152334642), 64'(-7686383409257), 64'(-4559778505553668), 64'(1089308448825112), 64'(171729321708043), 64'(-5460376320793), 64'(-5072342496187033), 64'(959328488094488), 64'(182520128106280), 64'(-3208428846785)},
		'{64'(-7789584925020678), 64'(-708887221199165), 64'(206702748225342), 64'(19845819841342), 64'(-7393588604643451), 64'(-873085743790196), 64'(189441643064668), 64'(21110141804838), 64'(-6918639246995094), 64'(-1024429359565484), 64'(170276674079431), 64'(22108944360992), 64'(-6371556198568998), 64'(-1161381434685658), 64'(149461551191327), 64'(22835111110925), 64'(-5759879607888814), 64'(-1282597644249583), 64'(127264837936296), 64'(23284800600436), 64'(-5091771080219080), 64'(-1386938313763298), 64'(103966594132105), 64'(23457435961283), 64'(-4375908801885863), 64'(-1473478185138064), 64'(79854941677743), 64'(23355656937656), 64'(-3621378440745346), 64'(-1541513537288910), 64'(55222594522994), 64'(22985235482840), 64'(-2837561156358186), 64'(-1590566623196775), 64'(30363393574260), 64'(22354956512905), 64'(-2034020064558654), 64'(-1620387416998168), 64'(5568886563148), 64'(21476465781009), 64'(-1220386496487468), 64'(-1630952695911038), 64'(-18875008286202), 64'(20364087183629), 64'(-406247372102900), 64'(-1622462512239951), 64'(-42691217575174), 64'(19034612125143), 64'(398965026813322), 64'(-1595334139989273), 64'(-65614571842050), 64'(17507063846682), 64'(1186079648425238), 64'(-1550193608429861), 64'(-87394675671863), 64'(15802439866299), 64'(1946288454422172), 64'(-1487864961015550), 64'(-107798558746634), 64'(13943435878177), 64'(2671242297735452), 64'(-1409357402058410), 64'(-126613080816760), 64'(11954154617207), 64'(3353139883456400), 64'(-1315850515302518), 64'(-143647066875011), 64'(9859803310540), 64'(3984808899006532), 64'(-1208677757771581), 64'(-158733152334649), 64'(7686383409256), 64'(4559778505553342), 64'(-1089308448825137), 64'(-171729321708049), 64'(5460376320792), 64'(5072342496186738), 64'(-959328488094511), 64'(-182520128106285), 64'(3208428846784)},
		'{64'(-20410122023596984), 64'(-1087203619517777), 64'(-261581401330405), 64'(-19688353631198), 64'(-19855845437227768), 64'(-1129165953014674), 64'(-260549776479662), 64'(-21497800075813), 64'(-19281639300793944), 64'(-1166937977762846), 64'(-258996978016206), 64'(-23185429430581), 64'(-18689575854732616), 64'(-1200612237457261), 64'(-256948048973282), 64'(-24752655664962), 64'(-18081679793730520), 64'(-1230286297560720), 64'(-254428064696757), 64'(-26201094598827), 64'(-17459925861202104), 64'(-1256062325165291), 64'(-251462077212791), 64'(-27532552007075), 64'(-16826236651983674), 64'(-1278046676369314), 64'(-248075061960339), 64'(-28749011807856), 64'(-16182480619338714), 64'(-1296349491750649), 64'(-244291866905447), 64'(-29852624356494), 64'(-15530470282089826), 64'(-1311084300475151), 64'(-240137164048391), 64'(-30845694866052), 64'(-14871960627433400), 64'(-1322367633538259), 64'(-235635403329143), 64'(-31730671974348), 64'(-14208647704754270), 64'(-1330318646597064), 64'(-230810768931151), 64'(-32510136476076), 64'(-13542167405539158), 64'(-1335058752810478), 64'(-225687137978284), 64'(-33186790237559), 64'(-12874094424288384), 64'(-1336711266066034), 64'(-220288041614798), 64'(-33763445310536), 64'(-12205941395145922), 64'(-1335401054933668), 64'(-214636628453457), 64'(-34243013260277), 64'(-11539158198806890), 64'(-1331254207649389), 64'(-208755630372409), 64'(-34628494722203), 64'(-10875131434119388), 64'(-1324397708395326), 64'(-202667330637182), 64'(-34922969200132), 64'(-10215184048673250), 64'(-1314959125107046), 64'(-196393534320064), 64'(-35129585118164), 64'(-9560575122561506), 64'(-1303066309004502), 64'(-189955540985356), 64'(-35251550137213), 64'(-8912499799410572), 64'(-1288847106009427), 64'(-183374119605357), 64'(-35292121746123), 64'(-8272089358702066), 64'(-1272429080179444), 64'(-176669485668604), 64'(-35254598136332)},
		'{64'(20410122023597112), 64'(1087203619517783), 64'(261581401330408), 64'(19688353631199), 64'(19855845437227944), 64'(1129165953014683), 64'(260549776479665), 64'(21497800075814), 64'(19281639300794168), 64'(1166937977762856), 64'(258996978016210), 64'(23185429430582), 64'(18689575854732880), 64'(1200612237457274), 64'(256948048973287), 64'(24752655664963), 64'(18081679793730820), 64'(1230286297560734), 64'(254428064696763), 64'(26201094598828), 64'(17459925861202444), 64'(1256062325165307), 64'(251462077212797), 64'(27532552007076), 64'(16826236651984046), 64'(1278046676369332), 64'(248075061960346), 64'(28749011807857), 64'(16182480619339120), 64'(1296349491750668), 64'(244291866905454), 64'(29852624356495), 64'(15530470282090264), 64'(1311084300475172), 64'(240137164048399), 64'(30845694866053), 64'(14871960627433864), 64'(1322367633538281), 64'(235635403329152), 64'(31730671974350), 64'(14208647704754760), 64'(1330318646597088), 64'(230810768931160), 64'(32510136476078), 64'(13542167405539672), 64'(1335058752810502), 64'(225687137978293), 64'(33186790237561), 64'(12874094424288920), 64'(1336711266066060), 64'(220288041614808), 64'(33763445310538), 64'(12205941395146478), 64'(1335401054933694), 64'(214636628453467), 64'(34243013260279), 64'(11539158198807466), 64'(1331254207649416), 64'(208755630372419), 64'(34628494722205), 64'(10875131434119980), 64'(1324397708395354), 64'(202667330637193), 64'(34922969200134), 64'(10215184048673856), 64'(1314959125107074), 64'(196393534320075), 64'(35129585118166), 64'(9560575122562122), 64'(1303066309004531), 64'(189955540985367), 64'(35251550137215), 64'(8912499799411199), 64'(1288847106009456), 64'(183374119605368), 64'(35292121746125), 64'(8272089358702702), 64'(1272429080179473), 64'(176669485668615), 64'(35254598136334)}};
	localparam logic signed[63:0] hf[0:1999] = {64'(7033096503296), 64'(-32897980416), 64'(-10967230464), 64'(63928604), 64'(7000245665792), 64'(-98394423296), 64'(-10337267712), 64'(188110032), 64'(6934845456384), 64'(-162997501952), 64'(-9086782464), 64'(301512896), 64'(6837488844800), 64'(-226124627968), 64'(-7233756672), 64'(397524544), 64'(6709056110592), 64'(-287210536960), 64'(-4804252672), 64'(470098240), 64'(6550703833088), 64'(-345713672192), 64'(-1831931776), 64'(513814560), 64'(6363853881344), 64'(-401122131968), 64'(1642511488), 64'(523933696), 64'(6150172966912), 64'(-452959338496), 64'(5571985920), 64'(496438560), 64'(5911558488064), 64'(-500788854784), 64'(9903706112), 64'(428068320), 64'(5650113888256), 64'(-544219168768), 64'(14579948544), 64'(316342016), 64'(5368126111744), 64'(-582907527168), 64'(19538849792), 64'(159572240), 64'(5068042010624), 64'(-616563212288), 64'(24715249664), 64'(-43130884), 64'(4752438460416), 64'(-644950327296), 64'(30041542656), 64'(-291865696), 64'(4423997194240), 64'(-667889827840), 64'(35448557568), 64'(-585954240), 64'(4085474918400), 64'(-685260537856), 64'(40866439168), 64'(-923966848), 64'(3739673690112), 64'(-697000263680), 64'(46225510400), 64'(-1303755136), 64'(3389412343808), 64'(-703105531904), 64'(51457126400), 64'(-1722493184), 64'(3037497131008), 64'(-703630671872), 64'(56494514176), 64'(-2176726784), 64'(2686692360192), 64'(-698686832640), 64'(61273546752), 64'(-2662427904), 64'(2339693658112), 64'(-688439820288), 64'(65733513216), 64'(-3175056896), 64'(1999099920384), 64'(-673107279872), 64'(69817778176), 64'(-3709628672), 64'(1667389456384), 64'(-652956008448), 64'(73474457600), 64'(-4260784384), 64'(1346895216640), 64'(-628297957376), 64'(76656959488), 64'(-4822863872), 64'(1039784017920), 64'(-599486234624), 64'(79324479488), 64'(-5389984768), 64'(748036685824), 64'(-566910648320), 64'(81442447360), 64'(-5956117504), 64'(473431015424), 64'(-530992660480), 64'(82982838272), 64'(-6515166720), 64'(217527091200), 64'(-492180406272), 64'(83924451328), 64'(-7061048320), 64'(-18344486912), 64'(-450943287296), 64'(84253073408), 64'(-7587765248), 64'(-233092038656), 64'(-407766368256), 64'(83961561088), 64'(-8089484800), 64'(-425869180928), 64'(-363144806400), 64'(83049857024), 64'(-8560607232), 64'(-596078428160), 64'(-317578280960), 64'(81524924416), 64'(-8995835904), 64'(-743372095488), 64'(-271565209600), 64'(79400542208), 64'(-9390236672), 64'(-867650306048), 64'(-225597456384), 64'(76697108480), 64'(-9739302912), 64'(-969056190464), 64'(-180154810368), 64'(73441320960), 64'(-10038998016), 64'(-1047968874496), 64'(-135700045824), 64'(69665783808), 64'(-10285808640), 64'(-1104993583104), 64'(-92673966080), 64'(65408569344), 64'(-10476781568), 64'(-1140949254144), 64'(-51490967552), 64'(60712722432), 64'(-10609551360), 64'(-1156854972416), 64'(-12534914048), 64'(55625695232), 64'(-10682369024), 64'(-1153913061376), 64'(23844581376), 64'(50198769664), 64'(-10694119424), 64'(-1133491388416), 64'(57335398400), 64'(44486422528), 64'(-10644324352), 64'(-1097103966208), 64'(87665672192), 64'(38545653760), 64'(-10533150720), 64'(-1046390308864), 64'(114606071808), 64'(32435316736), 64'(-10361399296), 64'(-983093477376), 64'(137971515392), 64'(26215440384), 64'(-10130492416), 64'(-909037731840), 64'(157622370304), 64'(19946518528), 64'(-9842454528), 64'(-826105724928), 64'(173465124864), 64'(13688829952), 64'(-9499883520), 64'(-736215171072), 64'(185452544000), 64'(7501764608), 64'(-9105917952), 64'(-641296105472), 64'(193583169536), 64'(1443165440), 64'(-8664196096), 64'(-543267749888), 64'(197900484608), 64'(-4431298048), 64'(-8178812416), 64'(-444016885760), 64'(198491455488), 64'(-10068722688), 64'(-7654265856), 64'(-345376227328), 64'(195484614656), 64'(-15419525120), 64'(-7095408640), 64'(-249104269312), 64'(189047783424), 64'(-20437946368), 64'(-6507388928), 64'(-156866412544), 64'(179385237504), 64'(-25082505216), 64'(-5895589888), 64'(-70217392128), 64'(166734675968), 64'(-29316399104), 64'(-5265568768), 64'(9414508544), 64'(151363747840), 64'(-33107843072), 64'(-4622995968), 64'(80741564416), 64'(133566259200), 64'(-36430344192), 64'(-3973589248), 64'(142628683776), 64'(113658347520), 64'(-39262916608), 64'(-3323052544), 64'(194103558144), 64'(91974221824), 64'(-41590218752), 64'(-2677014272), 64'(234364616704), 64'(68861943808), 64'(-43402641408), 64'(-2040966400), 64'(262786842624), 64'(44679032832), 64'(-44696309760), 64'(-1420208256), 64'(278925475840), 64'(19788113920), 64'(-45473042432), 64'(-819790720), 64'(282517438464), 64'(-5447470592), 64'(-45740224512), 64'(-244465792), 64'(273480531968), 64'(-30667960320), 64'(-45510623232), 64'(301360416), 64'(251910750208), 64'(-55521345536), 64'(-44802162688), 64'(813669824), 64'(218077265920), 64'(-79667380224), 64'(-43637624832), 64'(1288869760), 64'(172415664128), 64'(-102781378560), 64'(-42044309504), 64'(1723824640), 64'(115519225856), 64'(-124557795328), 64'(-40053633024), 64'(2115882240), 64'(48128520192), 64'(-144713433088), 64'(-37700722688), 64'(2462894336), 64'(-28880474112), 64'(-162990424064), 64'(-35023921152), 64'(2763230464), 64'(-114509742080), 64'(-179158859776), 64'(-32064319488), 64'(3015787008), 64'(-207653748736), 64'(-193018920960), 64'(-28865234944), 64'(3219988736), 64'(-307115032576), 64'(-204402835456), 64'(-25471664128), 64'(3375784960), 64'(-411620442112), 64'(-213176172544), 64'(-21929756672), 64'(3483641344), 64'(-519838269440), 64'(-219238973440), 64'(-18286260224), 64'(3544522240), 64'(-630395568128), 64'(-222526259200), 64'(-14587981824), 64'(3559872512), 64'(-741895634944), 64'(-223008227328), 64'(-10881244160), 64'(3531590144), 64'(-852935704576), 64'(-220690022400), 64'(-7211374080), 64'(3461996544), 64'(-962124054528), 64'(-215611097088), 64'(-3622200320), 64'(3353801728), 64'(-1068097273856), 64'(-207844130816), 64'(-155578656), 64'(3210066176), 64'(-1169536057344), 64'(-197493669888), 64'(3149049344), 64'(3034159104), 64'(-1265181130752), 64'(-184694308864), 64'(6255063040), 64'(2829713920), 64'(-1353847668736), 64'(-169608675328), 64'(9129030656), 64'(2600581376), 64'(-1434438467584), 64'(-152425005056), 64'(11741032448), 64'(2350781696), 64'(-1505956593664), 64'(-133354577920), 64'(14064936960), 64'(2084455552), 64'(-1567515475968), 64'(-112628752384), 64'(16078633984), 64'(1805813376), 64'(-1618349129728), 64'(-90496016384), 64'(17764208640), 64'(1519086592), 64'(-1657819234304), 64'(-67218747392), 64'(19108071424), 64'(1228478592), 64'(-1685421162496), 64'(-43069902848), 64'(20101029888), 64'(938116672), 64'(-1700789092352), 64'(-18329671680), 64'(20738314240), 64'(652006464), 64'(-1703698104320), 64'(6717959680), 64'(21019545600), 64'(373988160), 64'(-1694065885184), 64'(31788576768), 64'(20948656128), 64'(107695488), 64'(-1671951417344), 64'(56600698880), 64'(20533766144), 64'(-143481952), 64'(-1637553012736), 64'(80879017984), 64'(19787003904), 64'(-376432992), 64'(-1591204642816), 64'(104357543936), 64'(18724286464), 64'(-588355264), 64'(-1533370171392), 64'(126782562304), 64'(17365071872), 64'(-776781440), 64'(-1464636669952), 64'(147915423744), 64'(15732052992), 64'(-939601280), 64'(-1385706160128), 64'(167535099904), 64'(13850836992), 64'(-1075078784), 64'(-1297386569728), 64'(185440518144), 64'(11749591040), 64'(-1181864704), 64'(-1200580722688), 64'(201452535808), 64'(9458661376), 64'(-1259004928), 64'(-1096275197952), 64'(215415816192), 64'(7010174464), 64'(-1305943424), 64'(-985527877632), 64'(227200188416), 64'(4437632000), 64'(-1322520576), 64'(-869455364096), 64'(236701794304), 64'(1775485824), 64'(-1308967168), 64'(-749219348480), 64'(243843940352), 64'(-941283776), 64'(-1265894400), 64'(-626012913664), 64'(248577572864), 64'(-3677590016), 64'(-1194278144), 64'(-501046935552), 64'(250881425408), 64'(-6398656512), 64'(-1095440768), 64'(-375535730688), 64'(250761838592), 64'(-9070423040), 64'(-971028672), 64'(-250683834368), 64'(248252301312), 64'(-11659934720), 64'(-822986240), 64'(-127672295424), 64'(243412647936), 64'(-14135713792), 64'(-653526912), 64'(-7645917696), 64'(236328009728), 64'(-16468104192), 64'(-465101920), 64'(108299083776), 64'(227107389440), 64'(-18629595136), 64'(-260366176), 64'(219126661120), 64'(215882104832), 64'(-20595109888), 64'(-42143052), 64'(323871637504), 64'(202803920896), 64'(-22342254592), 64'(186612704), 64'(421649350656), 64'(188043018240), 64'(-23851552768), 64'(422852640), 64'(511664455680), 64'(171785748480), 64'(-25106614272), 64'(663472896), 64'(593218240512), 64'(154232242176), 64'(-26094284800), 64'(905352320), 64'(665715081216), 64'(135593918464), 64'(-26804754432), 64'(1145390336), 64'(728667193344), 64'(116090904576), 64'(-27231608832), 64'(1380543744), 64'(781698727936), 64'(95949373440), 64'(-27371864064), 64'(1607862400), 64'(824547606528), 64'(75398856704), 64'(-27225939968), 64'(1824522752), 64'(857067028480), 64'(54669598720), 64'(-26797602816), 64'(2027859968), 64'(879224750080), 64'(33989888000), 64'(-26093875200), 64'(2215397376), 64'(891101773824), 64'(13583513600), 64'(-25124898816), 64'(2384873216), 64'(892889333760), 64'(-6332733440), 64'(-23903772672), 64'(2534263552), 64'(884884701184), 64'(-25551407104), 64'(-22446352384), 64'(2661804288), 64'(867486269440), 64'(-43876618240), 64'(-20771020800), 64'(2766007296), 64'(841186934784), 64'(-61126078464), 64'(-18898444288), 64'(2845674240), 64'(806566887424), 64'(-77132947456), 64'(-16851289088), 64'(2899907328), 64'(764285681664), 64'(-91747483648), 64'(-14653930496), 64'(2928114688), 64'(715073060864), 64'(-104838455296), 64'(-12332148736), 64'(2930013696), 64'(659719585792), 64'(-116294311936), 64'(-9912799232), 64'(2905629696), 64'(599066345472), 64'(-126024146944), 64'(-7423496704), 64'(2855291904), 64'(533994668032), 64'(-133958361088), 64'(-4892274176), 64'(2779624704), 64'(465415241728), 64'(-140049088512), 64'(-2347257600), 64'(2679536640), 64'(394257203200), 64'(-144270393344), 64'(183660272), 64'(2556206336), 64'(321457225728), 64'(-146618138624), 64'(2673139712), 64'(2411064576), 64'(247948623872), 64'(-147109675008), 64'(5094700032), 64'(2245774336), 64'(174650785792), 64'(-145783259136), 64'(7423012352), 64'(2062207744), 64'(102458908672), 64'(-142697250816), 64'(9634170880), 64'(1862423296), 64'(32234213376), 64'(-137929080832), 64'(11705949184), 64'(1648637312), 64'(-35205341184), 64'(-131574038528), 64'(13618027520), 64'(1423197824), 64'(-99093577728), 64'(-123743797248), 64'(15352196096), 64'(1188554880), 64'(-158723964928), 64'(-114564939776), 64'(16892532736), 64'(947231424), 64'(-213456617472), 64'(-104177123328), 64'(18225549312), 64'(701792896), 64'(-262724354048), 64'(-92731334656), 64'(19340306432), 64'(454817568), 64'(-306037915648), 64'(-80387866624), 64'(20228497408), 64'(208866800), 64'(-342990127104), 64'(-67314339840), 64'(20884506624), 64'(-33544018), 64'(-373259010048), 64'(-53683642368), 64'(21305427968), 64'(-269973504), 64'(-396609880064), 64'(-39671808000), 64'(21491048448), 64'(-498081024), 64'(-412896460800), 64'(-25455941632), 64'(21443817472), 64'(-715651776), 64'(-422060851200), 64'(-11212149760), 64'(21168769024), 64'(-920620160), 64'(-424132542464), 64'(2886491648), 64'(20673421312), 64'(-1111091072), 64'(-419226353664), 64'(16671883264), 64'(19967651840), 64'(-1285358592), 64'(-407539548160), 64'(29982767104), 64'(19063545856), 64'(-1441922816), 64'(-389347966976), 64'(42666471424), 64'(17975222272), 64'(-1579503232), 64'(-365001244672), 64'(54580543488), 64'(16718628864), 64'(-1697049984), 64'(-334917435392), 64'(65594208256), 64'(15311344640), 64'(-1793752448), 64'(-299576754176), 64'(75589697536), 64'(13772339200), 64'(-1869043840), 64'(-259514777600), 64'(84463378432), 64'(12121732096), 64'(-1922604416), 64'(-215315218432), 64'(92126724096), 64'(10380551168), 64'(-1954360704), 64'(-167602061312), 64'(98507071488), 64'(8570467840), 64'(-1964482176), 64'(-117031575552), 64'(103548190720), 64'(6713540096), 64'(-1953375744), 64'(-64283930624), 64'(107210645504), 64'(4831954432), 64'(-1921676416), 64'(-10054776832), 64'(109471981568), 64'(2947766016), 64'(-1870237312), 64'(44953247744), 64'(110326685696), 64'(1082651264), 64'(-1800114816), 64'(100038934528), 64'(109785948160), 64'(-742337920), 64'(-1712554752), 64'(154510770176), 64'(107877253120), 64'(-2507003392), 64'(-1608973312), 64'(207694921728), 64'(104643788800), 64'(-4192218624), 64'(-1490939392), 64'(258942943232), 64'(100143644672), 64'(-5780130304), 64'(-1360152832), 64'(307638960128), 64'(94448910336), 64'(-7254341120), 64'(-1218423808), 64'(353206403072), 64'(87644585984), 64'(-8600073216), 64'(-1067649472), 64'(395114184704), 64'(79827378176), 64'(-9804311552), 64'(-909791232), 64'(432882253824), 64'(71104356352), 64'(-10855919616), 64'(-746850816), 64'(466086363136), 64'(61591547904), 64'(-11745739776), 64'(-580847104), 64'(494362230784), 64'(51412426752), 64'(-12466658304), 64'(-413792224), 64'(517408784384), 64'(40696356864), 64'(-13013656576), 64'(-247669072), 64'(534990848000), 64'(29576974336), 64'(-13383830528), 64'(-84408840), 64'(546940780544), 64'(18190557184), 64'(-13576387584), 64'(74130096), 64'(553159360512), 64'(6674405888), 64'(-13592614912), 64'(226182256), 64'(553615949824), 64'(-4834780672), 64'(-13435834368), 64'(370093632), 64'(548347740160), 64'(-16202491904), 64'(-13111324672), 64'(504338656), 64'(537458442240), 64'(-27297931264), 64'(-12626223104), 64'(627535488), 64'(521115828224), 64'(-37995479040), 64'(-11989416960), 64'(738459264), 64'(499548880896), 64'(-48176078848), 64'(-11211404288), 64'(836053504), 64'(473044221952), 64'(-57728499712), 64'(-10304146432), 64'(919438912), 64'(441941950464), 64'(-66550517760), 64'(-9280902144), 64'(987920768), 64'(406630694912), 64'(-74549952512), 64'(-8156052992), 64'(1040993088), 64'(367542566912), 64'(-81645584384), 64'(-6944914944), 64'(1078341504), 64'(325147328512), 64'(-87767891968), 64'(-5663543808), 64'(1099843200), 64'(279946461184), 64'(-92859727872), 64'(-4328539136), 64'(1105564672), 64'(232466825216), 64'(-96876699648), 64'(-2956838144), 64'(1095757824), 64'(183254220800), 64'(-99787579392), 64'(-1565513600), 64'(1070853440), 64'(132866760704), 64'(-101574352896), 64'(-171574784), 64'(1031453312), 64'(81868210176), 64'(-102232301568), 64'(1208231424), 64'(978319616), 64'(30821447680), 64'(-101769781248), 64'(2557609472), 64'(912363520), 64'(-19718068224), 64'(-100207943680), 64'(3860898560), 64'(834631680), 64'(-69208547328), 64'(-97580294144), 64'(5103242240), 64'(746291840), 64'(-117127929856), 64'(-93932068864), 64'(6270749696), 64'(648616768), 64'(-162979545088), 64'(-89319563264), 64'(7350639104), 64'(542967744), 64'(-206297481216), 64'(-83809280000), 64'(8331369472), 64'(430777056), 64'(-246651437056), 64'(-77476986880), 64'(9202753536), 64'(313529888), 64'(-283651080192), 64'(-70406725632), 64'(9956050944), 64'(192746128), 64'(-316949954560), 64'(-62689660928), 64'(10584052736), 64'(69961976), 64'(-346248708096), 64'(-54422949888), 64'(11081128960), 64'(-53288364), 64'(-371297878016), 64'(-45708509184), 64'(11443279872), 64'(-175490560), 64'(-391899774976), 64'(-36651757568), 64'(11668144128), 64'(-295167552), 64'(-407910121472), 64'(-27360344064), 64'(11755006976), 64'(-410896192), 64'(-419238739968), 64'(-17942872064), 64'(11704777728), 64'(-521323040), 64'(-425849716736), 64'(-8507630592), 64'(11519951872), 64'(-625179008), 64'(-427760877568), 64'(838650880), 64'(11204558848), 64'(-721292672), 64'(-425042903040), 64'(9992007680), 64'(10764085248), 64'(-808602688), 64'(-417817427968), 64'(18852395008), 64'(10205391872), 64'(-886167872), 64'(-406254944256), 64'(27324768256), 64'(9536608256), 64'(-953176704), 64'(-390571982848), 64'(35320111104), 64'(8767017984), 64'(-1008954368), 64'(-371027836928), 64'(42756349952), 64'(7906931200), 64'(-1052968640), 64'(-347921055744), 64'(49559191552), 64'(6967550976), 64'(-1084833536), 64'(-321585086464), 64'(55662837760), 64'(5960825344), 64'(-1104311424), 64'(-292384145408), 64'(61010624512), 64'(4899297280), 64'(-1111313664), 64'(-260708253696), 64'(65555509248), 64'(3795950592), 64'(-1105899136), 64'(-226968616960), 64'(69260451840), 64'(2664050688), 64'(-1088270976), 64'(-191592300544), 64'(72098676736), 64'(1516986752), 64'(-1058772032), 64'(-155017199616), 64'(74053804032), 64'(368114528), 64'(-1017878592), 64'(-117686788096), 64'(75119886336), 64'(-769398208), 64'(-966192896), 64'(-80044908544), 64'(75301273600), 64'(-1882721152), 64'(-904433792), 64'(-42530721792), 64'(74612400128), 64'(-2959504384), 64'(-833426688), 64'(-5573702144), 64'(73077473280), 64'(-3988013824), 64'(-754092160), 64'(30411114496), 64'(70729965568), 64'(-4957257216), 64'(-667433984), 64'(65027657728), 64'(67612160000), 64'(-5857098752), 64'(-574525888), 64'(97903050752), 64'(63774429184), 64'(-6678363136), 64'(-476498048), 64'(128691486720), 64'(59274575872), 64'(-7412924928), 64'(-374523168), 64'(157077749760), 64'(54177009664), 64'(-8053787136), 64'(-269802144), 64'(182780313600), 64'(48551907328), 64'(-8595142656), 64'(-163549664), 64'(205553975296), 64'(42474287104), 64'(-9032420352), 64'(-56980000), 64'(225192067072), 64'(36023083008), 64'(-9362321408), 64'(48707084), 64'(241528176640), 64'(29280149504), 64'(-9582834688), 64'(152339968), 64'(254437326848), 64'(22329272320), 64'(-9693236224), 64'(252788304), 64'(263836680192), 64'(15255162880), 64'(-9694081024), 64'(348975392), 64'(269685833728), 64'(8142476288), 64'(-9587174400), 64'(439889728), 64'(271986458624), 64'(1074818560), 64'(-9375527936), 64'(524595744), 64'(270781579264), 64'(-5866192896), 64'(-9063308288), 64'(602243328), 64'(266154344448), 64'(-12601840640), 64'(-8655766528), 64'(672076160), 64'(258226323456), 64'(-19057170432), 64'(-8159164928), 64'(733439296), 64'(247155507200), 64'(-25161789440), 64'(-7580680704), 64'(785784512), 64'(233133752320), 64'(-30850611200), 64'(-6928315392), 64'(828675456), 64'(216383995904), 64'(-36064505856), 64'(-6210783744), 64'(861790464), 64'(197157126144), 64'(-40750891008), 64'(-5437403136), 64'(884924608), 64'(175728607232), 64'(-44864233472), 64'(-4617976320), 64'(897990272), 64'(152394776576), 64'(-48366440448), 64'(-3762670080), 64'(901015872), 64'(127469125632), 64'(-51227189248), 64'(-2881891584), 64'(894144000), 64'(101278294016), 64'(-53424144384), 64'(-1986164096), 64'(877627648), 64'(74158080000), 64'(-54943068160), 64'(-1086004096), 64'(851825792), 64'(46449369088), 64'(-55777853440), 64'(-191799792), 64'(817197120), 64'(18494062592), 64'(-55930470400), 64'(686306496), 64'(774293504), 64'(-9368892416), 64'(-55410786304), 64'(1538531200), 64'(723751744), 64'(-36807413760), 64'(-54236319744), 64'(2355556864), 64'(666285184), 64'(-63500029952), 64'(-52431921152), 64'(3128631040), 64'(602673856), 64'(-89139437568), 64'(-50029350912), 64'(3849658368), 64'(533754816), 64'(-113435836416), 64'(-47066787840), 64'(4511283200), 64'(460411168), 64'(-136120008704), 64'(-43588292608), 64'(5106960896), 64'(383561312), 64'(-156946137088), 64'(-39643185152), 64'(5631021568), 64'(304147840), 64'(-175694184448), 64'(-35285385216), 64'(6078718976), 64'(223126112), 64'(-192172146688), 64'(-30572709888), 64'(6446269952), 64'(141453168), 64'(-206217691136), 64'(-25566150656), 64'(6730883584), 64'(60076656), 64'(-217699647488), 64'(-20329084928), 64'(6930774016), 64'(-20075964), 64'(-226518974464), 64'(-14926526464), 64'(7045166592), 64'(-98107728), 64'(-232609366016), 64'(-9424327680), 64'(7074288128), 64'(-173161984), 64'(-235937497088), 64'(-3888407296), 64'(7019345920), 64'(-244431584), 64'(-236502859776), 64'(1616015232), 64'(6882502144), 64'(-311167360), 64'(-234337206272), 64'(7025165824), 64'(6666826240), 64'(-372685728), 64'(-229503696896), 64'(12277432320), 64'(6376248320), 64'(-428375552), 64'(-222095589376), 64'(17314041856), 64'(6015498752), 64'(-477703744), 64'(-212234715136), 64'(22079696896), 64'(5590036992), 64'(-520220320), 64'(-200069513216), 64'(26523152384), 64'(5105980416), 64'(-555562048), 64'(-185772982272), 64'(30597754880), 64'(4570017280), 64'(-583455104), 64'(-169540141056), 64'(34261897216), 64'(3989324800), 64'(-603716864), 64'(-151585505280), 64'(37479415808), 64'(3371473408), 64'(-616256256), 64'(-132140228608), 64'(40219930624), 64'(2724335104), 64'(-621073344), 64'(-111449161728), 64'(42459090944), 64'(2055986048), 64'(-618257728), 64'(-89767772160), 64'(44178755584), 64'(1374610176), 64'(-607985920), 64'(-67359031296), 64'(45367111680), 64'(688401792), 64'(-590518080), 64'(-44490215424), 64'(46018699264), 64'(5471468), 64'(-566193024), 64'(-21429762048), 64'(46134370304), 64'(-666247424), 64'(-535423520), 64'(1555883136), 64'(45721169920), 64'(-1319086976), 64'(-498689888), 64'(24205301760), 64'(44792164352), 64'(-1945729536), 64'(-456533408), 64'(46265061376), 64'(43366166528), 64'(-2539286272), 64'(-409548928), 64'(67492519936), 64'(41467457536), 64'(-3093369600), 64'(-358377120), 64'(87658446848), 64'(39125377024), 64'(-3602159872), 64'(-303696256), 64'(106549485568), 64'(36373929984), 64'(-4060461568), 64'(-246213632), 64'(123970330624), 64'(33251299328), 64'(-4463754240), 64'(-186656976), 64'(139745705984), 64'(29799337984), 64'(-4808232448), 64'(-125765560), 64'(153722093568), 64'(26063024128), 64'(-5090839552), 64'(-64281496), 64'(165769084928), 64'(22089889792), 64'(-5309289472), 64'(-2941044), 64'(175780577280), 64'(17929424896), 64'(-5462078464), 64'(57533836), 64'(183675584512), 64'(13632480256), 64'(-5548493312), 64'(116443600), 64'(189398745088), 64'(9250644992), 64'(-5568603136), 64'(173118880), 64'(192920535040), 64'(4835645952), 64'(-5523246592), 64'(226927712), 64'(194237251584), 64'(438742560), 64'(-5414009344), 64'(277282272), 64'(193370537984), 64'(-3889856000), 64'(-5243192832), 64'(323644960), 64'(190366760960), 64'(-8101555712), 64'(-5013775360), 64'(365533728), 64'(185296093184), 64'(-12149912576), 64'(-4729367040), 64'(402526848), 64'(178251268096), 64'(-15991135232), 64'(-4394157056), 64'(434266688), 64'(169346187264), 64'(-19584544768), 64'(-4012854528), 64'(460462816), 64'(158714167296), 64'(-22892994560), 64'(-3590626816), 64'(480894272), 64'(146506186752), 64'(-25883242496), 64'(-3133030656), 64'(495411008), 64'(132888772608), 64'(-28526272512), 64'(-2645941760), 64'(503934304), 64'(118041862144), 64'(-30797553664), 64'(-2135481216), 64'(506456576), 64'(102156492800), 64'(-32677253120), 64'(-1607940736), 64'(503040352), 64'(85432393728), 64'(-34150387712), 64'(-1069706688), 64'(493816192), 64'(68075581440), 64'(-35206914048), 64'(-527184576), 64'(478980192), 64'(50295820288), 64'(-35841761280), 64'(13275691), 64'(458790528), 64'(32304191488), 64'(-36054810624), 64'(545452224), 64'(433563520), 64'(14310600704), 64'(-35850821632), 64'(1063321216), 64'(403668896), 64'(-3478606336), 64'(-35239272448), 64'(1561123456), 64'(369524608), 64'(-20862973952), 64'(-34234189824), 64'(2033426688), 64'(331591296), 64'(-37650149376), 64'(-32853913600), 64'(2475182848), 64'(290366144), 64'(-53657956352), 64'(-31120795648), 64'(2881780480), 64'(246376544), 64'(-68716351488), 64'(-29060892672), 64'(3249091072), 64'(200173424), 64'(-82669150208), 64'(-26703589376), 64'(3573507840), 64'(152324528), 64'(-95375622144), 64'(-24081211392), 64'(3851980032), 64'(103407576), 64'(-106711851008), 64'(-21228597248), 64'(4082038528), 64'(54003312), 64'(-116571865088), 64'(-18182653952), 64'(4261814272), 64'(4688806), 64'(-124868567040), 64'(-14981902336), 64'(4390051328), 64'(-43969216), 64'(-131534446592), 64'(-11665993728), 64'(4466109440), 64'(-91420760), 64'(-136521965568), 64'(-8275239936), 64'(4489962496), 64'(-137138640), 64'(-139803836416), 64'(-4850135552), 64'(4462188544), 64'(-180624272), 64'(-141372964864), 64'(-1430882688), 64'(4383951872), 64'(-221412864), 64'(-141242171392), 64'(1943064960), 64'(4256981760), 64'(-259078384), 64'(-139443732480), 64'(5233448448), 64'(4083541248), 64'(-293237696), 64'(-136028684288), 64'(8403623936), 64'(3866393344), 64'(-323554464), 64'(-131065856000), 64'(11418961920), 64'(3608760064), 64'(-349742080), 64'(-124640845824), 64'(14247211008), 64'(3314277632), 64'(-371566368), 64'(-116854710272), 64'(16858833920), 64'(2986947328), 64'(-388847200), 64'(-107822514176), 64'(19227299840), 64'(2631084288), 64'(-401459936), 64'(-97671798784), 64'(21329344512), 64'(2251260672), 64'(-409335712), 64'(-86540869632), 64'(23145181184), 64'(1852249216), 64'(-412461504), 64'(-74577018880), 64'(24658677760), 64'(1438965504), 64'(-410879232), 64'(-61934665728), 64'(25857468416), 64'(1016407424), 64'(-404684448), 64'(-48773451776), 64'(26733047808), 64'(589596736), 64'(-394024256), 64'(-35256303616), 64'(27280797696), 64'(163520480), 64'(-379094880), 64'(-21547479040), 64'(27499972608), 64'(-256926192), 64'(-360138432), 64'(-7810651136), 64'(27393648640), 64'(-666995136), 64'(-337439520), 64'(5792974336), 64'(26968619008), 64'(-1062137472), 64'(-311321088), 64'(19106494464), 64'(26235260928), 64'(-1438052992), 64'(-282140192), 64'(31979048960), 64'(25207339008), 64'(-1790736000), 64'(-250283168), 64'(44267466752), 64'(23901808640), 64'(-2116516096), 64'(-216160832), 64'(55837798400), 64'(22338547712), 64'(-2412095488), 64'(-180203184), 64'(66566709248), 64'(20540094464), 64'(-2674580480), 64'(-142854208), 64'(76342730752), 64'(18531325952), 64'(-2901509120), 64'(-104566496), 64'(85067358208), 64'(16339141632), 64'(-3090871296), 64'(-65795828), 64'(92655960064), 64'(13992113152), 64'(-3241124864), 64'(-26995910), 64'(99038543872), 64'(11520123904), 64'(-3351205888), 64'(11386859), 64'(104160296960), 64'(8954007552), 64'(-3420532224), 64'(48918428), 64'(107981996032), 64'(6325167616), 64'(-3449003264), 64'(85181896), 64'(110480179200), 64'(3665207808), 64'(-3436992256), 64'(119782032), 64'(111647170560), 64'(1005561408), 64'(-3385333760), 64'(152349504), 64'(111490867200), 64'(-1622868352), 64'(-3295307008), 64'(182544688), 64'(110034436096), 64'(-4190059008), 64'(-3168613632), 64'(210061120), 64'(107315757056), 64'(-6667201024), 64'(-3007350016), 64'(234628432), 64'(103386734592), 64'(-9027011584), 64'(-2813977088), 64'(256014944), 64'(98312503296), 64'(-11244024832), 64'(-2591285760), 64'(274029632), 64'(92170379264), 64'(-13294855168), 64'(-2342358784), 64'(288523648), 64'(85048827904), 64'(-15158435840), 64'(-2070530560), 64'(299391392), 64'(77046226944), 64'(-16816222208), 64'(-1779343616), 64'(306570976), 64'(68269547520), 64'(-18252363776), 64'(-1472505088), 64'(310044160), 64'(58832982016), 64'(-19453847552), 64'(-1153840384), 64'(309835904), 64'(48856506368), 64'(-20410593280), 64'(-827246976), 64'(306013216), 64'(38464389120), 64'(-21115523072), 64'(-496648352), 64'(298683904), 64'(27783663616), 64'(-21564604416), 64'(-165947968), 64'(287994368), 64'(16942639104), 64'(-21756829696), 64'(161015488), 64'(274127456), 64'(6069367296), 64'(-21694183424), 64'(480511552), 64'(257299680), 64'(-4709823488), 64'(-21381576704), 64'(788959168), 64'(237758064), 64'(-15271768064), 64'(-20826730496), 64'(1082965888), 64'(215776896), 64'(-25497839616), 64'(-20040044544), 64'(1359363712), 64'(191653968), 64'(-35275247616), 64'(-19034429440), 64'(1615242112), 64'(165706880), 64'(-44498239488), 64'(-17825124352), 64'(1847977472), 64'(138268864), 64'(-53069225984), 64'(-16429464576), 64'(2055258368), 64'(109684824), 64'(-60899762176), 64'(-14866663424), 64'(2235107584), 64'(80307000), 64'(-67911417856), 64'(-13157547008), 64'(2385898752), 64'(50490892), 64'(-74036527104), 64'(-11324291072), 64'(2506369792), 64'(20591002), 64'(-79218802688), 64'(-9390139392), 64'(2595631104), 64'(-9043209), 64'(-83413778432), 64'(-7379118592), 64'(2653169920), 64'(-38071296), 64'(-86589120512), 64'(-5315746304), 64'(2678849792), 64'(-66165620), 64'(-88724840448), 64'(-3224739072), 64'(2672905216), 64'(-93014920), 64'(-89813286912), 64'(-1130721792), 64'(2635934208), 64'(-118327656), 64'(-89859039232), 64'(942053824), 64'(2568883456), 64'(-141835040), 64'(-88878645248), 64'(2969985280), 64'(2473032960), 64'(-163293760), 64'(-86900252672), 64'(4930381312), 64'(2349974784), 64'(-182488384), 64'(-83963068416), 64'(6801708544), 64'(2201590016), 64'(-199233408), 64'(-80116711424), 64'(8563822592), 64'(2030020992), 64'(-213374832), 64'(-75420508160), 64'(10198177792), 64'(1837643904), 64'(-224791472), 64'(-69942599680), 64'(11688014848), 64'(1627035520), 64'(-233395808), 64'(-63759036416), 64'(13018524672), 64'(1400941312), 64'(-239134400), 64'(-56952745984), 64'(14176988160), 64'(1162240128), 64'(-241988000), 64'(-49612476416), 64'(15152887808), 64'(913908864), 64'(-241971088), 64'(-41831669760), 64'(15937992704), 64'(658986304), 64'(-239131280), 64'(-33707284480), 64'(16526415872), 64'(400536864), 64'(-233548080), 64'(-25338644480), 64'(16914642944), 64'(141614768), 64'(-225331520), 64'(-16826230784), 64'(17101535232), 64'(-114771248), 64'(-214620368), 64'(-8270504960), 64'(17088299008), 64'(-365691968), 64'(-201579968), 64'(229250672), 64'(16878435328), 64'(-608330368), 64'(-186399968), 64'(8576060928), 64'(16477662208), 64'(-840012160), 64'(-169291648), 64'(16676343808), 64'(15893807104), 64'(-1058234624), 64'(-150485136), 64'(24440932352), 64'(15136688128), 64'(-1260692480), 64'(-130226448), 64'(31786033152), 64'(14217958400), 64'(-1445301760), 64'(-108774312), 64'(38634110976), 64'(13150946304), 64'(-1610219392), 64'(-86397032), 64'(44914671616), 64'(11950475264), 64'(-1753861248), 64'(-63369172), 64'(50564964352), 64'(10632657920), 64'(-1874915968), 64'(-39968276), 64'(55530573824), 64'(9214700544), 64'(-1972355584), 64'(-16471616), 64'(59765919744), 64'(7714673664), 64'(-2045442560), 64'(6847026), 64'(63234625536), 64'(6151298560), 64'(-2093733376), 64'(29720462), 64'(65909788672), 64'(4543711744), 64'(-2117079296), 64'(51891092), 64'(67774132224), 64'(2911243008), 64'(-2115622528), 64'(73113720), 64'(68820041728), 64'(1273183616), 64'(-2089790208), 64'(93158192), 64'(69049499648), 64'(-351433280), 64'(-2040284416), 64'(111811808), 64'(68473896960), 64'(-1944049536), 64'(-1968069376), 64'(128881496), 64'(67113725952), 64'(-3486789120), 64'(-1874356352), 64'(144195728), 64'(64998219776), 64'(-4962652672), 64'(-1760584960), 64'(157606112), 64'(62164844544), 64'(-6355700736), 64'(-1628403200), 64'(168988784), 64'(58658750464), 64'(-7651218944), 64'(-1479644416), 64'(178245392), 64'(54532087808), 64'(-8835868672), 64'(-1316303360), 64'(185303792), 64'(49843318784), 64'(-9897820160), 64'(-1140510208), 64'(190118496), 64'(44656418816), 64'(-10826858496), 64'(-954503680), 64'(192670752), 64'(39040032768), 64'(-11614480384), 64'(-760603392), 64'(192968256), 64'(33066635264), 64'(-12253963264), 64'(-561181504), 64'(191044672), 64'(26811590656), 64'(-12740410368), 64'(-358634592), 64'(186958800), 64'(20352258048), 64'(-13070778368), 64'(-155355344), 64'(180793488), 64'(13767048192), 64'(-13243881472), 64'(46295076), 64'(172654240), 64'(7134508032), 64'(-13260374016), 64'(244013680), 64'(162667648), 64'(532402080), 64'(-13122712576), 64'(435581472), 64'(150979568), 64'(-5963171840), 64'(-12835095552), 64'(618887680), 64'(137753088), 64'(-12278635520), 64'(-12403388416), 64'(791952384), 64'(123166384), 64'(-18343737344), 64'(-11835023360), 64'(952947136), 64'(107410400), 64'(-24092315648), 64'(-11138892800), 64'(1100213760), 64'(90686408), 64'(-29462990848), 64'(-10325217280), 64'(1232280576), 64'(73203528), 64'(-34399793152), 64'(-9405405184), 64'(1347876480), 64'(55176152), 64'(-38852730880), 64'(-8391904768), 64'(1445942016), 64'(36821416), 64'(-42778251264), 64'(-7298036736), 64'(1525638272), 64'(18356602), 64'(-46139658240), 64'(-6137830912), 64'(1586352896), 64'(-3364), 64'(-48907403264), 64'(-4925849088), 64'(1627703296), 64'(-18048354), 64'(-51059314688), 64'(-3677007104), 64'(1649537408), 64'(-35575396), 64'(-52580737024), 64'(-2406398464), 64'(1651931392), 64'(-52390896), 64'(-53464559616), 64'(-1129114624), 64'(1635185152), 64'(-68312728), 64'(-53711183872), 64'(139928944), 64'(1599814784), 64'(-83172152), 64'(-53328396288), 64'(1386162304), 64'(1546543488), 64'(-96815528), 64'(-52331134976), 64'(2595524096), 64'(1476289152), 64'(-109105848), 64'(-50741219328), 64'(3754616064), 64'(1390150784), 64'(-119924056), 64'(-48586973184), 64'(4850846208), 64'(1289392896), 64'(-129170104), 64'(-45902774272), 64'(5872562688), 64'(1175427840), 64'(-136763808), 64'(-42728583168), 64'(6809170432), 64'(1049796992), 64'(-142645424), 64'(-39109353472), 64'(7651239424), 64'(914150976), 64'(-146776032), 64'(-35094458368), 64'(8390590464), 64'(770228544), 64'(-149137584), 64'(-30737025024), 64'(9020372992), 64'(619834944), 64'(-149732832), 64'(-26093264896), 64'(9535118336), 64'(464820192), 64'(-148584864), 64'(-21221765120), 64'(9930782720), 64'(307056544), 64'(-145736576), 64'(-16182777856), 64'(10204768256), 64'(148416656), 64'(-141249808), 64'(-11037487104), 64'(10355931136), 64'(-9248055), 64'(-135204288), 64'(-5847291392), 64'(10384567296), 64'(-164128624), 64'(-127696448), 64'(-673083584), 64'(10292387840), 64'(-314478656), 64'(-118838032), 64'(4425443328), 64'(10082473984), 64'(-458633504), 64'(-108754496), 64'(9390467072), 64'(9759219712), 64'(-595028224), 64'(-97583376), 64'(14166675456), 64'(9328256000), 64'(-722214016), 64'(-85472480), 64'(18701864960), 64'(8796367872), 64'(-838872960), 64'(-72578000), 64'(22947489792), 64'(8171397632), 64'(-943831040), 64'(-59062548), 64'(26859171840), 64'(7462130688), 64'(-1036069504), 64'(-45093212), 64'(30397132800), 64'(6678184448), 64'(-1114734080), 64'(-30839494), 64'(33526589440), 64'(5829879808), 64'(-1179141760), 64'(-16471352), 64'(36218060800), 64'(4928109056), 64'(-1228786048), 64'(-2157196), 64'(38447636480), 64'(3984203008), 64'(-1263340160), 64'(11938022), 64'(40197140480), 64'(3009790464), 64'(-1282657280), 64'(25654662), 64'(41454268416), 64'(2016659712), 64'(-1286769408), 64'(38840152), 64'(42212614144), 64'(1016618176), 64'(-1275884288), 64'(51350640), 64'(42471653376), 64'(21356334), 64'(-1250379776), 64'(63052516), 64'(42236645376), 64'(-957685888), 64'(-1210796416), 64'(73823768), 64'(41518489600), 64'(-1909447296), 64'(-1157828864), 64'(83555224), 64'(40333484032), 64'(-2823367424), 64'(-1092315392), 64'(92151592), 64'(38703067136), 64'(-3689500160), 64'(-1015224960), 64'(99532312), 64'(36653469696), 64'(-4498618368), 64'(-927644736), 64'(105632264), 64'(34215340032), 64'(-5242309120), 64'(-830765056), 64'(110402272), 64'(31423309824), 64'(-5913057792), 64'(-725863872), 64'(113809368), 64'(28315527168), 64'(-6504319488), 64'(-614290688), 64'(115836928), 64'(24933158912), 64'(-7010576896), 64'(-497449664), 64'(116484592), 64'(21319860224), 64'(-7427391488), 64'(-376782464), 64'(115767992), 64'(17521235968), 64'(-7751432704), 64'(-253750912), 64'(113718288), 64'(13584269312), 64'(-7980498432), 64'(-129819680), 64'(110381560), 64'(9556759552), 64'(-8113524224), 64'(-6439408), 64'(105818040), 64'(5486758400), 64'(-8150574080), 64'(114969968), 64'(100101136), 64'(1422006400), 64'(-8092821504), 64'(233035072), 64'(93316416), 64'(-2590614528), 64'(-7942518272), 64'(346444256), 64'(85560352), 64'(-6505608704), 64'(-7702948864), 64'(453961664), 64'(76939064), 64'(-10279368704), 64'(-7378376192), 64'(554440448), 64'(67566928), 64'(-13870651392), 64'(-6973975552), 64'(646834304), 64'(57565096), 64'(-17241012224), 64'(-6495759872), 64'(730208128), 64'(47059976), 64'(-20355205120), 64'(-5950494720), 64'(803746816), 64'(36181704), 64'(-23181537280), 64'(-5345609216), 64'(866762944), 64'(25062552), 64'(-25692176384), 64'(-4689098240), 64'(918702144), 64'(13835381), 64'(-27863408640), 64'(-3989420544), 64'(959147840), 64'(2632072), 64'(-29675841536), 64'(-3255392000), 64'(987823232), 64'(-8417969), 64'(-31114557440), 64'(-2496078848), 64'(1004592512), 64'(-19189274), 64'(-32169211904), 64'(-1720688896), 64'(1009460096), 64'(-29561700), 64'(-32834078720), 64'(-938460864), 64'(1002568000), 64'(-39421732), 64'(-33108035584), 64'(-158558640), 64'(984192000), 64'(-48663680), 64'(-32994498560), 64'(610034432), 64'(954736192), 64'(-57190776)};
	localparam logic signed[63:0] hb[0:1999] = {64'(7033096503296), 64'(32897980416), 64'(-10967230464), 64'(-63928604), 64'(7000245665792), 64'(98394423296), 64'(-10337267712), 64'(-188110032), 64'(6934845456384), 64'(162997501952), 64'(-9086782464), 64'(-301512896), 64'(6837488844800), 64'(226124627968), 64'(-7233756672), 64'(-397524544), 64'(6709056110592), 64'(287210536960), 64'(-4804252672), 64'(-470098240), 64'(6550703833088), 64'(345713672192), 64'(-1831931776), 64'(-513814560), 64'(6363853881344), 64'(401122131968), 64'(1642511488), 64'(-523933696), 64'(6150172966912), 64'(452959338496), 64'(5571985920), 64'(-496438560), 64'(5911558488064), 64'(500788854784), 64'(9903706112), 64'(-428068320), 64'(5650113888256), 64'(544219168768), 64'(14579948544), 64'(-316342016), 64'(5368126111744), 64'(582907527168), 64'(19538849792), 64'(-159572240), 64'(5068042010624), 64'(616563212288), 64'(24715249664), 64'(43130884), 64'(4752438460416), 64'(644950327296), 64'(30041542656), 64'(291865696), 64'(4423997194240), 64'(667889827840), 64'(35448557568), 64'(585954240), 64'(4085474918400), 64'(685260537856), 64'(40866439168), 64'(923966848), 64'(3739673690112), 64'(697000263680), 64'(46225510400), 64'(1303755136), 64'(3389412343808), 64'(703105531904), 64'(51457126400), 64'(1722493184), 64'(3037497131008), 64'(703630671872), 64'(56494514176), 64'(2176726784), 64'(2686692360192), 64'(698686832640), 64'(61273546752), 64'(2662427904), 64'(2339693658112), 64'(688439820288), 64'(65733513216), 64'(3175056896), 64'(1999099920384), 64'(673107279872), 64'(69817778176), 64'(3709628672), 64'(1667389456384), 64'(652956008448), 64'(73474457600), 64'(4260784384), 64'(1346895216640), 64'(628297957376), 64'(76656959488), 64'(4822863872), 64'(1039784017920), 64'(599486234624), 64'(79324479488), 64'(5389984768), 64'(748036685824), 64'(566910648320), 64'(81442447360), 64'(5956117504), 64'(473431015424), 64'(530992660480), 64'(82982838272), 64'(6515166720), 64'(217527091200), 64'(492180406272), 64'(83924451328), 64'(7061048320), 64'(-18344486912), 64'(450943287296), 64'(84253073408), 64'(7587765248), 64'(-233092038656), 64'(407766368256), 64'(83961561088), 64'(8089484800), 64'(-425869180928), 64'(363144806400), 64'(83049857024), 64'(8560607232), 64'(-596078428160), 64'(317578280960), 64'(81524924416), 64'(8995835904), 64'(-743372095488), 64'(271565209600), 64'(79400542208), 64'(9390236672), 64'(-867650306048), 64'(225597456384), 64'(76697108480), 64'(9739302912), 64'(-969056190464), 64'(180154810368), 64'(73441320960), 64'(10038998016), 64'(-1047968874496), 64'(135700045824), 64'(69665783808), 64'(10285808640), 64'(-1104993583104), 64'(92673966080), 64'(65408569344), 64'(10476781568), 64'(-1140949254144), 64'(51490967552), 64'(60712722432), 64'(10609551360), 64'(-1156854972416), 64'(12534914048), 64'(55625695232), 64'(10682369024), 64'(-1153913061376), 64'(-23844581376), 64'(50198769664), 64'(10694119424), 64'(-1133491388416), 64'(-57335398400), 64'(44486422528), 64'(10644324352), 64'(-1097103966208), 64'(-87665672192), 64'(38545653760), 64'(10533150720), 64'(-1046390308864), 64'(-114606071808), 64'(32435316736), 64'(10361399296), 64'(-983093477376), 64'(-137971515392), 64'(26215440384), 64'(10130492416), 64'(-909037731840), 64'(-157622370304), 64'(19946518528), 64'(9842454528), 64'(-826105724928), 64'(-173465124864), 64'(13688829952), 64'(9499883520), 64'(-736215171072), 64'(-185452544000), 64'(7501764608), 64'(9105917952), 64'(-641296105472), 64'(-193583169536), 64'(1443165440), 64'(8664196096), 64'(-543267749888), 64'(-197900484608), 64'(-4431298048), 64'(8178812416), 64'(-444016885760), 64'(-198491455488), 64'(-10068722688), 64'(7654265856), 64'(-345376227328), 64'(-195484614656), 64'(-15419525120), 64'(7095408640), 64'(-249104269312), 64'(-189047783424), 64'(-20437946368), 64'(6507388928), 64'(-156866412544), 64'(-179385237504), 64'(-25082505216), 64'(5895589888), 64'(-70217392128), 64'(-166734675968), 64'(-29316399104), 64'(5265568768), 64'(9414508544), 64'(-151363747840), 64'(-33107843072), 64'(4622995968), 64'(80741564416), 64'(-133566259200), 64'(-36430344192), 64'(3973589248), 64'(142628683776), 64'(-113658347520), 64'(-39262916608), 64'(3323052544), 64'(194103558144), 64'(-91974221824), 64'(-41590218752), 64'(2677014272), 64'(234364616704), 64'(-68861943808), 64'(-43402641408), 64'(2040966400), 64'(262786842624), 64'(-44679032832), 64'(-44696309760), 64'(1420208256), 64'(278925475840), 64'(-19788113920), 64'(-45473042432), 64'(819790720), 64'(282517438464), 64'(5447470592), 64'(-45740224512), 64'(244465792), 64'(273480531968), 64'(30667960320), 64'(-45510623232), 64'(-301360416), 64'(251910750208), 64'(55521345536), 64'(-44802162688), 64'(-813669824), 64'(218077265920), 64'(79667380224), 64'(-43637624832), 64'(-1288869760), 64'(172415664128), 64'(102781378560), 64'(-42044309504), 64'(-1723824640), 64'(115519225856), 64'(124557795328), 64'(-40053633024), 64'(-2115882240), 64'(48128520192), 64'(144713433088), 64'(-37700722688), 64'(-2462894336), 64'(-28880474112), 64'(162990424064), 64'(-35023921152), 64'(-2763230464), 64'(-114509742080), 64'(179158859776), 64'(-32064319488), 64'(-3015787008), 64'(-207653748736), 64'(193018920960), 64'(-28865234944), 64'(-3219988736), 64'(-307115032576), 64'(204402835456), 64'(-25471664128), 64'(-3375784960), 64'(-411620442112), 64'(213176172544), 64'(-21929756672), 64'(-3483641344), 64'(-519838269440), 64'(219238973440), 64'(-18286260224), 64'(-3544522240), 64'(-630395568128), 64'(222526259200), 64'(-14587981824), 64'(-3559872512), 64'(-741895634944), 64'(223008227328), 64'(-10881244160), 64'(-3531590144), 64'(-852935704576), 64'(220690022400), 64'(-7211374080), 64'(-3461996544), 64'(-962124054528), 64'(215611097088), 64'(-3622200320), 64'(-3353801728), 64'(-1068097273856), 64'(207844130816), 64'(-155578656), 64'(-3210066176), 64'(-1169536057344), 64'(197493669888), 64'(3149049344), 64'(-3034159104), 64'(-1265181130752), 64'(184694308864), 64'(6255063040), 64'(-2829713920), 64'(-1353847668736), 64'(169608675328), 64'(9129030656), 64'(-2600581376), 64'(-1434438467584), 64'(152425005056), 64'(11741032448), 64'(-2350781696), 64'(-1505956593664), 64'(133354577920), 64'(14064936960), 64'(-2084455552), 64'(-1567515475968), 64'(112628752384), 64'(16078633984), 64'(-1805813376), 64'(-1618349129728), 64'(90496016384), 64'(17764208640), 64'(-1519086592), 64'(-1657819234304), 64'(67218747392), 64'(19108071424), 64'(-1228478592), 64'(-1685421162496), 64'(43069902848), 64'(20101029888), 64'(-938116672), 64'(-1700789092352), 64'(18329671680), 64'(20738314240), 64'(-652006464), 64'(-1703698104320), 64'(-6717959680), 64'(21019545600), 64'(-373988160), 64'(-1694065885184), 64'(-31788576768), 64'(20948656128), 64'(-107695488), 64'(-1671951417344), 64'(-56600698880), 64'(20533766144), 64'(143481952), 64'(-1637553012736), 64'(-80879017984), 64'(19787003904), 64'(376432992), 64'(-1591204642816), 64'(-104357543936), 64'(18724286464), 64'(588355264), 64'(-1533370171392), 64'(-126782562304), 64'(17365071872), 64'(776781440), 64'(-1464636669952), 64'(-147915423744), 64'(15732052992), 64'(939601280), 64'(-1385706160128), 64'(-167535099904), 64'(13850836992), 64'(1075078784), 64'(-1297386569728), 64'(-185440518144), 64'(11749591040), 64'(1181864704), 64'(-1200580722688), 64'(-201452535808), 64'(9458661376), 64'(1259004928), 64'(-1096275197952), 64'(-215415816192), 64'(7010174464), 64'(1305943424), 64'(-985527877632), 64'(-227200188416), 64'(4437632000), 64'(1322520576), 64'(-869455364096), 64'(-236701794304), 64'(1775485824), 64'(1308967168), 64'(-749219348480), 64'(-243843940352), 64'(-941283776), 64'(1265894400), 64'(-626012913664), 64'(-248577572864), 64'(-3677590016), 64'(1194278144), 64'(-501046935552), 64'(-250881425408), 64'(-6398656512), 64'(1095440768), 64'(-375535730688), 64'(-250761838592), 64'(-9070423040), 64'(971028672), 64'(-250683834368), 64'(-248252301312), 64'(-11659934720), 64'(822986240), 64'(-127672295424), 64'(-243412647936), 64'(-14135713792), 64'(653526912), 64'(-7645917696), 64'(-236328009728), 64'(-16468104192), 64'(465101920), 64'(108299083776), 64'(-227107389440), 64'(-18629595136), 64'(260366176), 64'(219126661120), 64'(-215882104832), 64'(-20595109888), 64'(42143052), 64'(323871637504), 64'(-202803920896), 64'(-22342254592), 64'(-186612704), 64'(421649350656), 64'(-188043018240), 64'(-23851552768), 64'(-422852640), 64'(511664455680), 64'(-171785748480), 64'(-25106614272), 64'(-663472896), 64'(593218240512), 64'(-154232242176), 64'(-26094284800), 64'(-905352320), 64'(665715081216), 64'(-135593918464), 64'(-26804754432), 64'(-1145390336), 64'(728667193344), 64'(-116090904576), 64'(-27231608832), 64'(-1380543744), 64'(781698727936), 64'(-95949373440), 64'(-27371864064), 64'(-1607862400), 64'(824547606528), 64'(-75398856704), 64'(-27225939968), 64'(-1824522752), 64'(857067028480), 64'(-54669598720), 64'(-26797602816), 64'(-2027859968), 64'(879224750080), 64'(-33989888000), 64'(-26093875200), 64'(-2215397376), 64'(891101773824), 64'(-13583513600), 64'(-25124898816), 64'(-2384873216), 64'(892889333760), 64'(6332733440), 64'(-23903772672), 64'(-2534263552), 64'(884884701184), 64'(25551407104), 64'(-22446352384), 64'(-2661804288), 64'(867486269440), 64'(43876618240), 64'(-20771020800), 64'(-2766007296), 64'(841186934784), 64'(61126078464), 64'(-18898444288), 64'(-2845674240), 64'(806566887424), 64'(77132947456), 64'(-16851289088), 64'(-2899907328), 64'(764285681664), 64'(91747483648), 64'(-14653930496), 64'(-2928114688), 64'(715073060864), 64'(104838455296), 64'(-12332148736), 64'(-2930013696), 64'(659719585792), 64'(116294311936), 64'(-9912799232), 64'(-2905629696), 64'(599066345472), 64'(126024146944), 64'(-7423496704), 64'(-2855291904), 64'(533994668032), 64'(133958361088), 64'(-4892274176), 64'(-2779624704), 64'(465415241728), 64'(140049088512), 64'(-2347257600), 64'(-2679536640), 64'(394257203200), 64'(144270393344), 64'(183660272), 64'(-2556206336), 64'(321457225728), 64'(146618138624), 64'(2673139712), 64'(-2411064576), 64'(247948623872), 64'(147109675008), 64'(5094700032), 64'(-2245774336), 64'(174650785792), 64'(145783259136), 64'(7423012352), 64'(-2062207744), 64'(102458908672), 64'(142697250816), 64'(9634170880), 64'(-1862423296), 64'(32234213376), 64'(137929080832), 64'(11705949184), 64'(-1648637312), 64'(-35205341184), 64'(131574038528), 64'(13618027520), 64'(-1423197824), 64'(-99093577728), 64'(123743797248), 64'(15352196096), 64'(-1188554880), 64'(-158723964928), 64'(114564939776), 64'(16892532736), 64'(-947231424), 64'(-213456617472), 64'(104177123328), 64'(18225549312), 64'(-701792896), 64'(-262724354048), 64'(92731334656), 64'(19340306432), 64'(-454817568), 64'(-306037915648), 64'(80387866624), 64'(20228497408), 64'(-208866800), 64'(-342990127104), 64'(67314339840), 64'(20884506624), 64'(33544018), 64'(-373259010048), 64'(53683642368), 64'(21305427968), 64'(269973504), 64'(-396609880064), 64'(39671808000), 64'(21491048448), 64'(498081024), 64'(-412896460800), 64'(25455941632), 64'(21443817472), 64'(715651776), 64'(-422060851200), 64'(11212149760), 64'(21168769024), 64'(920620160), 64'(-424132542464), 64'(-2886491648), 64'(20673421312), 64'(1111091072), 64'(-419226353664), 64'(-16671883264), 64'(19967651840), 64'(1285358592), 64'(-407539548160), 64'(-29982767104), 64'(19063545856), 64'(1441922816), 64'(-389347966976), 64'(-42666471424), 64'(17975222272), 64'(1579503232), 64'(-365001244672), 64'(-54580543488), 64'(16718628864), 64'(1697049984), 64'(-334917435392), 64'(-65594208256), 64'(15311344640), 64'(1793752448), 64'(-299576754176), 64'(-75589697536), 64'(13772339200), 64'(1869043840), 64'(-259514777600), 64'(-84463378432), 64'(12121732096), 64'(1922604416), 64'(-215315218432), 64'(-92126724096), 64'(10380551168), 64'(1954360704), 64'(-167602061312), 64'(-98507071488), 64'(8570467840), 64'(1964482176), 64'(-117031575552), 64'(-103548190720), 64'(6713540096), 64'(1953375744), 64'(-64283930624), 64'(-107210645504), 64'(4831954432), 64'(1921676416), 64'(-10054776832), 64'(-109471981568), 64'(2947766016), 64'(1870237312), 64'(44953247744), 64'(-110326685696), 64'(1082651264), 64'(1800114816), 64'(100038934528), 64'(-109785948160), 64'(-742337920), 64'(1712554752), 64'(154510770176), 64'(-107877253120), 64'(-2507003392), 64'(1608973312), 64'(207694921728), 64'(-104643788800), 64'(-4192218624), 64'(1490939392), 64'(258942943232), 64'(-100143644672), 64'(-5780130304), 64'(1360152832), 64'(307638960128), 64'(-94448910336), 64'(-7254341120), 64'(1218423808), 64'(353206403072), 64'(-87644585984), 64'(-8600073216), 64'(1067649472), 64'(395114184704), 64'(-79827378176), 64'(-9804311552), 64'(909791232), 64'(432882253824), 64'(-71104356352), 64'(-10855919616), 64'(746850816), 64'(466086363136), 64'(-61591547904), 64'(-11745739776), 64'(580847104), 64'(494362230784), 64'(-51412426752), 64'(-12466658304), 64'(413792224), 64'(517408784384), 64'(-40696356864), 64'(-13013656576), 64'(247669072), 64'(534990848000), 64'(-29576974336), 64'(-13383830528), 64'(84408840), 64'(546940780544), 64'(-18190557184), 64'(-13576387584), 64'(-74130096), 64'(553159360512), 64'(-6674405888), 64'(-13592614912), 64'(-226182256), 64'(553615949824), 64'(4834780672), 64'(-13435834368), 64'(-370093632), 64'(548347740160), 64'(16202491904), 64'(-13111324672), 64'(-504338656), 64'(537458442240), 64'(27297931264), 64'(-12626223104), 64'(-627535488), 64'(521115828224), 64'(37995479040), 64'(-11989416960), 64'(-738459264), 64'(499548880896), 64'(48176078848), 64'(-11211404288), 64'(-836053504), 64'(473044221952), 64'(57728499712), 64'(-10304146432), 64'(-919438912), 64'(441941950464), 64'(66550517760), 64'(-9280902144), 64'(-987920768), 64'(406630694912), 64'(74549952512), 64'(-8156052992), 64'(-1040993088), 64'(367542566912), 64'(81645584384), 64'(-6944914944), 64'(-1078341504), 64'(325147328512), 64'(87767891968), 64'(-5663543808), 64'(-1099843200), 64'(279946461184), 64'(92859727872), 64'(-4328539136), 64'(-1105564672), 64'(232466825216), 64'(96876699648), 64'(-2956838144), 64'(-1095757824), 64'(183254220800), 64'(99787579392), 64'(-1565513600), 64'(-1070853440), 64'(132866760704), 64'(101574352896), 64'(-171574784), 64'(-1031453312), 64'(81868210176), 64'(102232301568), 64'(1208231424), 64'(-978319616), 64'(30821447680), 64'(101769781248), 64'(2557609472), 64'(-912363520), 64'(-19718068224), 64'(100207943680), 64'(3860898560), 64'(-834631680), 64'(-69208547328), 64'(97580294144), 64'(5103242240), 64'(-746291840), 64'(-117127929856), 64'(93932068864), 64'(6270749696), 64'(-648616768), 64'(-162979545088), 64'(89319563264), 64'(7350639104), 64'(-542967744), 64'(-206297481216), 64'(83809280000), 64'(8331369472), 64'(-430777056), 64'(-246651437056), 64'(77476986880), 64'(9202753536), 64'(-313529888), 64'(-283651080192), 64'(70406725632), 64'(9956050944), 64'(-192746128), 64'(-316949954560), 64'(62689660928), 64'(10584052736), 64'(-69961976), 64'(-346248708096), 64'(54422949888), 64'(11081128960), 64'(53288364), 64'(-371297878016), 64'(45708509184), 64'(11443279872), 64'(175490560), 64'(-391899774976), 64'(36651757568), 64'(11668144128), 64'(295167552), 64'(-407910121472), 64'(27360344064), 64'(11755006976), 64'(410896192), 64'(-419238739968), 64'(17942872064), 64'(11704777728), 64'(521323040), 64'(-425849716736), 64'(8507630592), 64'(11519951872), 64'(625179008), 64'(-427760877568), 64'(-838650880), 64'(11204558848), 64'(721292672), 64'(-425042903040), 64'(-9992007680), 64'(10764085248), 64'(808602688), 64'(-417817427968), 64'(-18852395008), 64'(10205391872), 64'(886167872), 64'(-406254944256), 64'(-27324768256), 64'(9536608256), 64'(953176704), 64'(-390571982848), 64'(-35320111104), 64'(8767017984), 64'(1008954368), 64'(-371027836928), 64'(-42756349952), 64'(7906931200), 64'(1052968640), 64'(-347921055744), 64'(-49559191552), 64'(6967550976), 64'(1084833536), 64'(-321585086464), 64'(-55662837760), 64'(5960825344), 64'(1104311424), 64'(-292384145408), 64'(-61010624512), 64'(4899297280), 64'(1111313664), 64'(-260708253696), 64'(-65555509248), 64'(3795950592), 64'(1105899136), 64'(-226968616960), 64'(-69260451840), 64'(2664050688), 64'(1088270976), 64'(-191592300544), 64'(-72098676736), 64'(1516986752), 64'(1058772032), 64'(-155017199616), 64'(-74053804032), 64'(368114528), 64'(1017878592), 64'(-117686788096), 64'(-75119886336), 64'(-769398208), 64'(966192896), 64'(-80044908544), 64'(-75301273600), 64'(-1882721152), 64'(904433792), 64'(-42530721792), 64'(-74612400128), 64'(-2959504384), 64'(833426688), 64'(-5573702144), 64'(-73077473280), 64'(-3988013824), 64'(754092160), 64'(30411114496), 64'(-70729965568), 64'(-4957257216), 64'(667433984), 64'(65027657728), 64'(-67612160000), 64'(-5857098752), 64'(574525888), 64'(97903050752), 64'(-63774429184), 64'(-6678363136), 64'(476498048), 64'(128691486720), 64'(-59274575872), 64'(-7412924928), 64'(374523168), 64'(157077749760), 64'(-54177009664), 64'(-8053787136), 64'(269802144), 64'(182780313600), 64'(-48551907328), 64'(-8595142656), 64'(163549664), 64'(205553975296), 64'(-42474287104), 64'(-9032420352), 64'(56980000), 64'(225192067072), 64'(-36023083008), 64'(-9362321408), 64'(-48707084), 64'(241528176640), 64'(-29280149504), 64'(-9582834688), 64'(-152339968), 64'(254437326848), 64'(-22329272320), 64'(-9693236224), 64'(-252788304), 64'(263836680192), 64'(-15255162880), 64'(-9694081024), 64'(-348975392), 64'(269685833728), 64'(-8142476288), 64'(-9587174400), 64'(-439889728), 64'(271986458624), 64'(-1074818560), 64'(-9375527936), 64'(-524595744), 64'(270781579264), 64'(5866192896), 64'(-9063308288), 64'(-602243328), 64'(266154344448), 64'(12601840640), 64'(-8655766528), 64'(-672076160), 64'(258226323456), 64'(19057170432), 64'(-8159164928), 64'(-733439296), 64'(247155507200), 64'(25161789440), 64'(-7580680704), 64'(-785784512), 64'(233133752320), 64'(30850611200), 64'(-6928315392), 64'(-828675456), 64'(216383995904), 64'(36064505856), 64'(-6210783744), 64'(-861790464), 64'(197157126144), 64'(40750891008), 64'(-5437403136), 64'(-884924608), 64'(175728607232), 64'(44864233472), 64'(-4617976320), 64'(-897990272), 64'(152394776576), 64'(48366440448), 64'(-3762670080), 64'(-901015872), 64'(127469125632), 64'(51227189248), 64'(-2881891584), 64'(-894144000), 64'(101278294016), 64'(53424144384), 64'(-1986164096), 64'(-877627648), 64'(74158080000), 64'(54943068160), 64'(-1086004096), 64'(-851825792), 64'(46449369088), 64'(55777853440), 64'(-191799792), 64'(-817197120), 64'(18494062592), 64'(55930470400), 64'(686306496), 64'(-774293504), 64'(-9368892416), 64'(55410786304), 64'(1538531200), 64'(-723751744), 64'(-36807413760), 64'(54236319744), 64'(2355556864), 64'(-666285184), 64'(-63500029952), 64'(52431921152), 64'(3128631040), 64'(-602673856), 64'(-89139437568), 64'(50029350912), 64'(3849658368), 64'(-533754816), 64'(-113435836416), 64'(47066787840), 64'(4511283200), 64'(-460411168), 64'(-136120008704), 64'(43588292608), 64'(5106960896), 64'(-383561312), 64'(-156946137088), 64'(39643185152), 64'(5631021568), 64'(-304147840), 64'(-175694184448), 64'(35285385216), 64'(6078718976), 64'(-223126112), 64'(-192172146688), 64'(30572709888), 64'(6446269952), 64'(-141453168), 64'(-206217691136), 64'(25566150656), 64'(6730883584), 64'(-60076656), 64'(-217699647488), 64'(20329084928), 64'(6930774016), 64'(20075964), 64'(-226518974464), 64'(14926526464), 64'(7045166592), 64'(98107728), 64'(-232609366016), 64'(9424327680), 64'(7074288128), 64'(173161984), 64'(-235937497088), 64'(3888407296), 64'(7019345920), 64'(244431584), 64'(-236502859776), 64'(-1616015232), 64'(6882502144), 64'(311167360), 64'(-234337206272), 64'(-7025165824), 64'(6666826240), 64'(372685728), 64'(-229503696896), 64'(-12277432320), 64'(6376248320), 64'(428375552), 64'(-222095589376), 64'(-17314041856), 64'(6015498752), 64'(477703744), 64'(-212234715136), 64'(-22079696896), 64'(5590036992), 64'(520220320), 64'(-200069513216), 64'(-26523152384), 64'(5105980416), 64'(555562048), 64'(-185772982272), 64'(-30597754880), 64'(4570017280), 64'(583455104), 64'(-169540141056), 64'(-34261897216), 64'(3989324800), 64'(603716864), 64'(-151585505280), 64'(-37479415808), 64'(3371473408), 64'(616256256), 64'(-132140228608), 64'(-40219930624), 64'(2724335104), 64'(621073344), 64'(-111449161728), 64'(-42459090944), 64'(2055986048), 64'(618257728), 64'(-89767772160), 64'(-44178755584), 64'(1374610176), 64'(607985920), 64'(-67359031296), 64'(-45367111680), 64'(688401792), 64'(590518080), 64'(-44490215424), 64'(-46018699264), 64'(5471468), 64'(566193024), 64'(-21429762048), 64'(-46134370304), 64'(-666247424), 64'(535423520), 64'(1555883136), 64'(-45721169920), 64'(-1319086976), 64'(498689888), 64'(24205301760), 64'(-44792164352), 64'(-1945729536), 64'(456533408), 64'(46265061376), 64'(-43366166528), 64'(-2539286272), 64'(409548928), 64'(67492519936), 64'(-41467457536), 64'(-3093369600), 64'(358377120), 64'(87658446848), 64'(-39125377024), 64'(-3602159872), 64'(303696256), 64'(106549485568), 64'(-36373929984), 64'(-4060461568), 64'(246213632), 64'(123970330624), 64'(-33251299328), 64'(-4463754240), 64'(186656976), 64'(139745705984), 64'(-29799337984), 64'(-4808232448), 64'(125765560), 64'(153722093568), 64'(-26063024128), 64'(-5090839552), 64'(64281496), 64'(165769084928), 64'(-22089889792), 64'(-5309289472), 64'(2941044), 64'(175780577280), 64'(-17929424896), 64'(-5462078464), 64'(-57533836), 64'(183675584512), 64'(-13632480256), 64'(-5548493312), 64'(-116443600), 64'(189398745088), 64'(-9250644992), 64'(-5568603136), 64'(-173118880), 64'(192920535040), 64'(-4835645952), 64'(-5523246592), 64'(-226927712), 64'(194237251584), 64'(-438742560), 64'(-5414009344), 64'(-277282272), 64'(193370537984), 64'(3889856000), 64'(-5243192832), 64'(-323644960), 64'(190366760960), 64'(8101555712), 64'(-5013775360), 64'(-365533728), 64'(185296093184), 64'(12149912576), 64'(-4729367040), 64'(-402526848), 64'(178251268096), 64'(15991135232), 64'(-4394157056), 64'(-434266688), 64'(169346187264), 64'(19584544768), 64'(-4012854528), 64'(-460462816), 64'(158714167296), 64'(22892994560), 64'(-3590626816), 64'(-480894272), 64'(146506186752), 64'(25883242496), 64'(-3133030656), 64'(-495411008), 64'(132888772608), 64'(28526272512), 64'(-2645941760), 64'(-503934304), 64'(118041862144), 64'(30797553664), 64'(-2135481216), 64'(-506456576), 64'(102156492800), 64'(32677253120), 64'(-1607940736), 64'(-503040352), 64'(85432393728), 64'(34150387712), 64'(-1069706688), 64'(-493816192), 64'(68075581440), 64'(35206914048), 64'(-527184576), 64'(-478980192), 64'(50295820288), 64'(35841761280), 64'(13275691), 64'(-458790528), 64'(32304191488), 64'(36054810624), 64'(545452224), 64'(-433563520), 64'(14310600704), 64'(35850821632), 64'(1063321216), 64'(-403668896), 64'(-3478606336), 64'(35239272448), 64'(1561123456), 64'(-369524608), 64'(-20862973952), 64'(34234189824), 64'(2033426688), 64'(-331591296), 64'(-37650149376), 64'(32853913600), 64'(2475182848), 64'(-290366144), 64'(-53657956352), 64'(31120795648), 64'(2881780480), 64'(-246376544), 64'(-68716351488), 64'(29060892672), 64'(3249091072), 64'(-200173424), 64'(-82669150208), 64'(26703589376), 64'(3573507840), 64'(-152324528), 64'(-95375622144), 64'(24081211392), 64'(3851980032), 64'(-103407576), 64'(-106711851008), 64'(21228597248), 64'(4082038528), 64'(-54003312), 64'(-116571865088), 64'(18182653952), 64'(4261814272), 64'(-4688806), 64'(-124868567040), 64'(14981902336), 64'(4390051328), 64'(43969216), 64'(-131534446592), 64'(11665993728), 64'(4466109440), 64'(91420760), 64'(-136521965568), 64'(8275239936), 64'(4489962496), 64'(137138640), 64'(-139803836416), 64'(4850135552), 64'(4462188544), 64'(180624272), 64'(-141372964864), 64'(1430882688), 64'(4383951872), 64'(221412864), 64'(-141242171392), 64'(-1943064960), 64'(4256981760), 64'(259078384), 64'(-139443732480), 64'(-5233448448), 64'(4083541248), 64'(293237696), 64'(-136028684288), 64'(-8403623936), 64'(3866393344), 64'(323554464), 64'(-131065856000), 64'(-11418961920), 64'(3608760064), 64'(349742080), 64'(-124640845824), 64'(-14247211008), 64'(3314277632), 64'(371566368), 64'(-116854710272), 64'(-16858833920), 64'(2986947328), 64'(388847200), 64'(-107822514176), 64'(-19227299840), 64'(2631084288), 64'(401459936), 64'(-97671798784), 64'(-21329344512), 64'(2251260672), 64'(409335712), 64'(-86540869632), 64'(-23145181184), 64'(1852249216), 64'(412461504), 64'(-74577018880), 64'(-24658677760), 64'(1438965504), 64'(410879232), 64'(-61934665728), 64'(-25857468416), 64'(1016407424), 64'(404684448), 64'(-48773451776), 64'(-26733047808), 64'(589596736), 64'(394024256), 64'(-35256303616), 64'(-27280797696), 64'(163520480), 64'(379094880), 64'(-21547479040), 64'(-27499972608), 64'(-256926192), 64'(360138432), 64'(-7810651136), 64'(-27393648640), 64'(-666995136), 64'(337439520), 64'(5792974336), 64'(-26968619008), 64'(-1062137472), 64'(311321088), 64'(19106494464), 64'(-26235260928), 64'(-1438052992), 64'(282140192), 64'(31979048960), 64'(-25207339008), 64'(-1790736000), 64'(250283168), 64'(44267466752), 64'(-23901808640), 64'(-2116516096), 64'(216160832), 64'(55837798400), 64'(-22338547712), 64'(-2412095488), 64'(180203184), 64'(66566709248), 64'(-20540094464), 64'(-2674580480), 64'(142854208), 64'(76342730752), 64'(-18531325952), 64'(-2901509120), 64'(104566496), 64'(85067358208), 64'(-16339141632), 64'(-3090871296), 64'(65795828), 64'(92655960064), 64'(-13992113152), 64'(-3241124864), 64'(26995910), 64'(99038543872), 64'(-11520123904), 64'(-3351205888), 64'(-11386859), 64'(104160296960), 64'(-8954007552), 64'(-3420532224), 64'(-48918428), 64'(107981996032), 64'(-6325167616), 64'(-3449003264), 64'(-85181896), 64'(110480179200), 64'(-3665207808), 64'(-3436992256), 64'(-119782032), 64'(111647170560), 64'(-1005561408), 64'(-3385333760), 64'(-152349504), 64'(111490867200), 64'(1622868352), 64'(-3295307008), 64'(-182544688), 64'(110034436096), 64'(4190059008), 64'(-3168613632), 64'(-210061120), 64'(107315757056), 64'(6667201024), 64'(-3007350016), 64'(-234628432), 64'(103386734592), 64'(9027011584), 64'(-2813977088), 64'(-256014944), 64'(98312503296), 64'(11244024832), 64'(-2591285760), 64'(-274029632), 64'(92170379264), 64'(13294855168), 64'(-2342358784), 64'(-288523648), 64'(85048827904), 64'(15158435840), 64'(-2070530560), 64'(-299391392), 64'(77046226944), 64'(16816222208), 64'(-1779343616), 64'(-306570976), 64'(68269547520), 64'(18252363776), 64'(-1472505088), 64'(-310044160), 64'(58832982016), 64'(19453847552), 64'(-1153840384), 64'(-309835904), 64'(48856506368), 64'(20410593280), 64'(-827246976), 64'(-306013216), 64'(38464389120), 64'(21115523072), 64'(-496648352), 64'(-298683904), 64'(27783663616), 64'(21564604416), 64'(-165947968), 64'(-287994368), 64'(16942639104), 64'(21756829696), 64'(161015488), 64'(-274127456), 64'(6069367296), 64'(21694183424), 64'(480511552), 64'(-257299680), 64'(-4709823488), 64'(21381576704), 64'(788959168), 64'(-237758064), 64'(-15271768064), 64'(20826730496), 64'(1082965888), 64'(-215776896), 64'(-25497839616), 64'(20040044544), 64'(1359363712), 64'(-191653968), 64'(-35275247616), 64'(19034429440), 64'(1615242112), 64'(-165706880), 64'(-44498239488), 64'(17825124352), 64'(1847977472), 64'(-138268864), 64'(-53069225984), 64'(16429464576), 64'(2055258368), 64'(-109684824), 64'(-60899762176), 64'(14866663424), 64'(2235107584), 64'(-80307000), 64'(-67911417856), 64'(13157547008), 64'(2385898752), 64'(-50490892), 64'(-74036527104), 64'(11324291072), 64'(2506369792), 64'(-20591002), 64'(-79218802688), 64'(9390139392), 64'(2595631104), 64'(9043209), 64'(-83413778432), 64'(7379118592), 64'(2653169920), 64'(38071296), 64'(-86589120512), 64'(5315746304), 64'(2678849792), 64'(66165620), 64'(-88724840448), 64'(3224739072), 64'(2672905216), 64'(93014920), 64'(-89813286912), 64'(1130721792), 64'(2635934208), 64'(118327656), 64'(-89859039232), 64'(-942053824), 64'(2568883456), 64'(141835040), 64'(-88878645248), 64'(-2969985280), 64'(2473032960), 64'(163293760), 64'(-86900252672), 64'(-4930381312), 64'(2349974784), 64'(182488384), 64'(-83963068416), 64'(-6801708544), 64'(2201590016), 64'(199233408), 64'(-80116711424), 64'(-8563822592), 64'(2030020992), 64'(213374832), 64'(-75420508160), 64'(-10198177792), 64'(1837643904), 64'(224791472), 64'(-69942599680), 64'(-11688014848), 64'(1627035520), 64'(233395808), 64'(-63759036416), 64'(-13018524672), 64'(1400941312), 64'(239134400), 64'(-56952745984), 64'(-14176988160), 64'(1162240128), 64'(241988000), 64'(-49612476416), 64'(-15152887808), 64'(913908864), 64'(241971088), 64'(-41831669760), 64'(-15937992704), 64'(658986304), 64'(239131280), 64'(-33707284480), 64'(-16526415872), 64'(400536864), 64'(233548080), 64'(-25338644480), 64'(-16914642944), 64'(141614768), 64'(225331520), 64'(-16826230784), 64'(-17101535232), 64'(-114771248), 64'(214620368), 64'(-8270504960), 64'(-17088299008), 64'(-365691968), 64'(201579968), 64'(229250672), 64'(-16878435328), 64'(-608330368), 64'(186399968), 64'(8576060928), 64'(-16477662208), 64'(-840012160), 64'(169291648), 64'(16676343808), 64'(-15893807104), 64'(-1058234624), 64'(150485136), 64'(24440932352), 64'(-15136688128), 64'(-1260692480), 64'(130226448), 64'(31786033152), 64'(-14217958400), 64'(-1445301760), 64'(108774312), 64'(38634110976), 64'(-13150946304), 64'(-1610219392), 64'(86397032), 64'(44914671616), 64'(-11950475264), 64'(-1753861248), 64'(63369172), 64'(50564964352), 64'(-10632657920), 64'(-1874915968), 64'(39968276), 64'(55530573824), 64'(-9214700544), 64'(-1972355584), 64'(16471616), 64'(59765919744), 64'(-7714673664), 64'(-2045442560), 64'(-6847026), 64'(63234625536), 64'(-6151298560), 64'(-2093733376), 64'(-29720462), 64'(65909788672), 64'(-4543711744), 64'(-2117079296), 64'(-51891092), 64'(67774132224), 64'(-2911243008), 64'(-2115622528), 64'(-73113720), 64'(68820041728), 64'(-1273183616), 64'(-2089790208), 64'(-93158192), 64'(69049499648), 64'(351433280), 64'(-2040284416), 64'(-111811808), 64'(68473896960), 64'(1944049536), 64'(-1968069376), 64'(-128881496), 64'(67113725952), 64'(3486789120), 64'(-1874356352), 64'(-144195728), 64'(64998219776), 64'(4962652672), 64'(-1760584960), 64'(-157606112), 64'(62164844544), 64'(6355700736), 64'(-1628403200), 64'(-168988784), 64'(58658750464), 64'(7651218944), 64'(-1479644416), 64'(-178245392), 64'(54532087808), 64'(8835868672), 64'(-1316303360), 64'(-185303792), 64'(49843318784), 64'(9897820160), 64'(-1140510208), 64'(-190118496), 64'(44656418816), 64'(10826858496), 64'(-954503680), 64'(-192670752), 64'(39040032768), 64'(11614480384), 64'(-760603392), 64'(-192968256), 64'(33066635264), 64'(12253963264), 64'(-561181504), 64'(-191044672), 64'(26811590656), 64'(12740410368), 64'(-358634592), 64'(-186958800), 64'(20352258048), 64'(13070778368), 64'(-155355344), 64'(-180793488), 64'(13767048192), 64'(13243881472), 64'(46295076), 64'(-172654240), 64'(7134508032), 64'(13260374016), 64'(244013680), 64'(-162667648), 64'(532402080), 64'(13122712576), 64'(435581472), 64'(-150979568), 64'(-5963171840), 64'(12835095552), 64'(618887680), 64'(-137753088), 64'(-12278635520), 64'(12403388416), 64'(791952384), 64'(-123166384), 64'(-18343737344), 64'(11835023360), 64'(952947136), 64'(-107410400), 64'(-24092315648), 64'(11138892800), 64'(1100213760), 64'(-90686408), 64'(-29462990848), 64'(10325217280), 64'(1232280576), 64'(-73203528), 64'(-34399793152), 64'(9405405184), 64'(1347876480), 64'(-55176152), 64'(-38852730880), 64'(8391904768), 64'(1445942016), 64'(-36821416), 64'(-42778251264), 64'(7298036736), 64'(1525638272), 64'(-18356602), 64'(-46139658240), 64'(6137830912), 64'(1586352896), 64'(3364), 64'(-48907403264), 64'(4925849088), 64'(1627703296), 64'(18048354), 64'(-51059314688), 64'(3677007104), 64'(1649537408), 64'(35575396), 64'(-52580737024), 64'(2406398464), 64'(1651931392), 64'(52390896), 64'(-53464559616), 64'(1129114624), 64'(1635185152), 64'(68312728), 64'(-53711183872), 64'(-139928944), 64'(1599814784), 64'(83172152), 64'(-53328396288), 64'(-1386162304), 64'(1546543488), 64'(96815528), 64'(-52331134976), 64'(-2595524096), 64'(1476289152), 64'(109105848), 64'(-50741219328), 64'(-3754616064), 64'(1390150784), 64'(119924056), 64'(-48586973184), 64'(-4850846208), 64'(1289392896), 64'(129170104), 64'(-45902774272), 64'(-5872562688), 64'(1175427840), 64'(136763808), 64'(-42728583168), 64'(-6809170432), 64'(1049796992), 64'(142645424), 64'(-39109353472), 64'(-7651239424), 64'(914150976), 64'(146776032), 64'(-35094458368), 64'(-8390590464), 64'(770228544), 64'(149137584), 64'(-30737025024), 64'(-9020372992), 64'(619834944), 64'(149732832), 64'(-26093264896), 64'(-9535118336), 64'(464820192), 64'(148584864), 64'(-21221765120), 64'(-9930782720), 64'(307056544), 64'(145736576), 64'(-16182777856), 64'(-10204768256), 64'(148416656), 64'(141249808), 64'(-11037487104), 64'(-10355931136), 64'(-9248055), 64'(135204288), 64'(-5847291392), 64'(-10384567296), 64'(-164128624), 64'(127696448), 64'(-673083584), 64'(-10292387840), 64'(-314478656), 64'(118838032), 64'(4425443328), 64'(-10082473984), 64'(-458633504), 64'(108754496), 64'(9390467072), 64'(-9759219712), 64'(-595028224), 64'(97583376), 64'(14166675456), 64'(-9328256000), 64'(-722214016), 64'(85472480), 64'(18701864960), 64'(-8796367872), 64'(-838872960), 64'(72578000), 64'(22947489792), 64'(-8171397632), 64'(-943831040), 64'(59062548), 64'(26859171840), 64'(-7462130688), 64'(-1036069504), 64'(45093212), 64'(30397132800), 64'(-6678184448), 64'(-1114734080), 64'(30839494), 64'(33526589440), 64'(-5829879808), 64'(-1179141760), 64'(16471352), 64'(36218060800), 64'(-4928109056), 64'(-1228786048), 64'(2157196), 64'(38447636480), 64'(-3984203008), 64'(-1263340160), 64'(-11938022), 64'(40197140480), 64'(-3009790464), 64'(-1282657280), 64'(-25654662), 64'(41454268416), 64'(-2016659712), 64'(-1286769408), 64'(-38840152), 64'(42212614144), 64'(-1016618176), 64'(-1275884288), 64'(-51350640), 64'(42471653376), 64'(-21356334), 64'(-1250379776), 64'(-63052516), 64'(42236645376), 64'(957685888), 64'(-1210796416), 64'(-73823768), 64'(41518489600), 64'(1909447296), 64'(-1157828864), 64'(-83555224), 64'(40333484032), 64'(2823367424), 64'(-1092315392), 64'(-92151592), 64'(38703067136), 64'(3689500160), 64'(-1015224960), 64'(-99532312), 64'(36653469696), 64'(4498618368), 64'(-927644736), 64'(-105632264), 64'(34215340032), 64'(5242309120), 64'(-830765056), 64'(-110402272), 64'(31423309824), 64'(5913057792), 64'(-725863872), 64'(-113809368), 64'(28315527168), 64'(6504319488), 64'(-614290688), 64'(-115836928), 64'(24933158912), 64'(7010576896), 64'(-497449664), 64'(-116484592), 64'(21319860224), 64'(7427391488), 64'(-376782464), 64'(-115767992), 64'(17521235968), 64'(7751432704), 64'(-253750912), 64'(-113718288), 64'(13584269312), 64'(7980498432), 64'(-129819680), 64'(-110381560), 64'(9556759552), 64'(8113524224), 64'(-6439408), 64'(-105818040), 64'(5486758400), 64'(8150574080), 64'(114969968), 64'(-100101136), 64'(1422006400), 64'(8092821504), 64'(233035072), 64'(-93316416), 64'(-2590614528), 64'(7942518272), 64'(346444256), 64'(-85560352), 64'(-6505608704), 64'(7702948864), 64'(453961664), 64'(-76939064), 64'(-10279368704), 64'(7378376192), 64'(554440448), 64'(-67566928), 64'(-13870651392), 64'(6973975552), 64'(646834304), 64'(-57565096), 64'(-17241012224), 64'(6495759872), 64'(730208128), 64'(-47059976), 64'(-20355205120), 64'(5950494720), 64'(803746816), 64'(-36181704), 64'(-23181537280), 64'(5345609216), 64'(866762944), 64'(-25062552), 64'(-25692176384), 64'(4689098240), 64'(918702144), 64'(-13835381), 64'(-27863408640), 64'(3989420544), 64'(959147840), 64'(-2632072), 64'(-29675841536), 64'(3255392000), 64'(987823232), 64'(8417969), 64'(-31114557440), 64'(2496078848), 64'(1004592512), 64'(19189274), 64'(-32169211904), 64'(1720688896), 64'(1009460096), 64'(29561700), 64'(-32834078720), 64'(938460864), 64'(1002568000), 64'(39421732), 64'(-33108035584), 64'(158558640), 64'(984192000), 64'(48663680), 64'(-32994498560), 64'(-610034432), 64'(954736192), 64'(57190776)};
endpackage
`endif
