`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam N = 4;
	localparam M = 4;
	localparam real Lfr[0:3] = {0.98900646, 0.98900646, 0.97591347, 0.97591347};
	localparam real Lfi[0:3] = {0.04798661, -0.04798661, 0.019232517, -0.019232517};
	localparam real Lbr[0:3] = {0.98900646, 0.98900646, 0.97591347, 0.97591347};
	localparam real Lbi[0:3] = {0.04798661, -0.04798661, 0.019232517, -0.019232517};
	localparam real Wfr[0:3] = {1.32158975e-05, 1.32158975e-05, -3.9246156e-06, -3.9246156e-06};
	localparam real Wfi[0:3] = {5.4198574e-07, -5.4198574e-07, -7.5876746e-06, 7.5876746e-06};
	localparam real Wbr[0:3] = {1.32158975e-05, 1.32158975e-05, 3.9246156e-06, 3.9246156e-06};
	localparam real Wbi[0:3] = {5.4198574e-07, -5.4198574e-07, 7.5876746e-06, -7.5876746e-06};
	localparam real Ffr[0:3][0:99] = '{
		'{183.25674, 17.803015, -1.9955642, 0.02115994, 191.84448, 16.545134, -2.006414, 0.027916582, 199.79929, 15.271762, -2.0121887, 0.034473382, 207.11423, 13.98629, -2.0129735, 0.040818363, 213.78412, 12.69207, -2.0088646, 0.046940286, 219.80539, 11.392408, -1.9999676, 0.05282868, 225.17615, 10.090563, -1.9863975, 0.058473844, 229.89612, 8.78973, -1.9682786, 0.06386685, 233.96657, 7.493044, -1.945744, 0.068999566, 237.39035, 6.2035656, -1.9189346, 0.073864646, 240.17183, 4.924279, -1.8879989, 0.07845553, 242.31682, 3.6580853, -1.8530928, 0.08276646, 243.83257, 2.4077973, -1.8143785, 0.086792454, 244.7277, 1.1761336, -1.7720243, 0.090529345, 245.01224, -0.03428483, -1.7262039, 0.093973726, 244.69739, -1.2209402, -1.6770965, 0.09712297, 243.79565, -2.3814216, -1.6248852, 0.09997521, 242.32071, -3.5134282, -1.5697573, 0.10252937, 240.28734, -4.614774, -1.5119035, 0.10478506, 237.71138, -5.683389, -1.4515173, 0.10674267, 234.60973, -6.7173247, -1.3887947, 0.10840329, 231.00014, -7.714753, -1.3239331, 0.109768696, 226.90134, -8.673971, -1.2571319, 0.110841356, 222.33281, -9.593401, -1.1885909, 0.111624405, 217.3148, -10.471594, -1.11851, 0.1121216},
		'{183.25674, 17.803015, -1.9955642, 0.02115994, 191.84448, 16.545134, -2.006414, 0.027916582, 199.79929, 15.271762, -2.0121887, 0.034473382, 207.11423, 13.98629, -2.0129735, 0.040818363, 213.78412, 12.69207, -2.0088646, 0.046940286, 219.80539, 11.392408, -1.9999676, 0.05282868, 225.17615, 10.090563, -1.9863975, 0.058473844, 229.89612, 8.78973, -1.9682786, 0.06386685, 233.96657, 7.493044, -1.945744, 0.068999566, 237.39035, 6.2035656, -1.9189346, 0.073864646, 240.17183, 4.924279, -1.8879989, 0.07845553, 242.31682, 3.6580853, -1.8530928, 0.08276646, 243.83257, 2.4077973, -1.8143785, 0.086792454, 244.7277, 1.1761336, -1.7720243, 0.090529345, 245.01224, -0.03428483, -1.7262039, 0.093973726, 244.69739, -1.2209402, -1.6770965, 0.09712297, 243.79565, -2.3814216, -1.6248852, 0.09997521, 242.32071, -3.5134282, -1.5697573, 0.10252937, 240.28734, -4.614774, -1.5119035, 0.10478506, 237.71138, -5.683389, -1.4515173, 0.10674267, 234.60973, -6.7173247, -1.3887947, 0.10840329, 231.00014, -7.714753, -1.3239331, 0.109768696, 226.90134, -8.673971, -1.2571319, 0.110841356, 222.33281, -9.593401, -1.1885909, 0.111624405, 217.3148, -10.471594, -1.11851, 0.1121216},
		'{-182.00656, -17.691608, 1.9211302, -0.2637629, -190.55325, -16.50202, 1.8158827, -0.2539327, -198.51532, -15.352927, 1.7138801, -0.2443255, -205.9128, -14.243513, 1.615066, -0.23493986, -212.7653, -13.172956, 1.5193839, -0.22577423, -219.09207, -12.14044, 1.4267766, -0.21682692, -224.91194, -11.145147, 1.3371872, -0.20809613, -230.24329, -10.186268, 1.2505579, -0.19957995, -235.10413, -9.262992, 1.1668315, -0.19127631, -239.51207, -8.374516, 1.0859503, -0.18318307, -243.48431, -7.520039, 1.0078568, -0.17529799, -247.03764, -6.6987696, 0.93249375, -0.16761872, -250.18848, -5.909919, 0.85980356, -0.16014284, -252.95282, -5.1527047, 0.7897292, -0.15286785, -255.34631, -4.4263535, 0.7222136, -0.14579117, -257.3842, -3.7300978, 0.6572003, -0.13891017, -259.0813, -3.0631773, 0.5946326, -0.13222215, -260.45212, -2.4248407, 0.5344547, -0.12572433, -261.51077, -1.8143445, 0.47661078, -0.11941391, -262.27097, -1.2309542, 0.42104563, -0.11328804, -262.74612, -0.67394376, 0.36770442, -0.10734382, -262.9492, -0.14259684, 0.3165328, -0.10157833, -262.89285, 0.3637938, 0.26747695, -0.095988594, -262.58945, 0.84592545, 0.22048353, -0.09057163, -262.05087, 1.3044858, 0.17549983, -0.08532442},
		'{-182.00656, -17.691608, 1.9211302, -0.2637629, -190.55325, -16.50202, 1.8158827, -0.2539327, -198.51532, -15.352927, 1.7138801, -0.2443255, -205.9128, -14.243513, 1.615066, -0.23493986, -212.7653, -13.172956, 1.5193839, -0.22577423, -219.09207, -12.14044, 1.4267766, -0.21682692, -224.91194, -11.145147, 1.3371872, -0.20809613, -230.24329, -10.186268, 1.2505579, -0.19957995, -235.10413, -9.262992, 1.1668315, -0.19127631, -239.51207, -8.374516, 1.0859503, -0.18318307, -243.48431, -7.520039, 1.0078568, -0.17529799, -247.03764, -6.6987696, 0.93249375, -0.16761872, -250.18848, -5.909919, 0.85980356, -0.16014284, -252.95282, -5.1527047, 0.7897292, -0.15286785, -255.34631, -4.4263535, 0.7222136, -0.14579117, -257.3842, -3.7300978, 0.6572003, -0.13891017, -259.0813, -3.0631773, 0.5946326, -0.13222215, -260.45212, -2.4248407, 0.5344547, -0.12572433, -261.51077, -1.8143445, 0.47661078, -0.11941391, -262.27097, -1.2309542, 0.42104563, -0.11328804, -262.74612, -0.67394376, 0.36770442, -0.10734382, -262.9492, -0.14259684, 0.3165328, -0.10157833, -262.89285, 0.3637938, 0.26747695, -0.095988594, -262.58945, 0.84592545, 0.22048353, -0.09057163, -262.05087, 1.3044858, 0.17549983, -0.08532442}};
	localparam real Ffi[0:3][0:99] = '{
		'{-220.94467, 22.134588, 0.68327236, -0.14565031, -209.72185, 22.745558, 0.58000046, -0.14303371, -198.2103, 23.28945, 0.4773432, -0.14012164, -186.44359, 23.766256, 0.3755374, -0.13692695, -174.4552, 24.176136, 0.27481315, -0.1334629, -162.27855, 24.519405, 0.17539336, -0.12974317, -149.94682, 24.796534, 0.0774935, -0.12578177, -137.49294, 25.008144, -0.018678905, -0.12159303, -124.94948, 25.155006, -0.11292458, -0.11719154, -112.34858, 25.23803, -0.20505281, -0.11259214, -99.72192, 25.258263, -0.29488173, -0.10780984, -87.100586, 25.216887, -0.3822386, -0.10285982, -74.51508, 25.115202, -0.4669601, -0.09775735, -61.9952, 24.954641, -0.54889244, -0.09251777, -49.570004, 24.73674, -0.62789166, -0.08715648, -37.267746, 24.463152, -0.70382357, -0.08168884, -25.115845, 24.135626, -0.77656424, -0.0761302, -13.140806, 23.756014, -0.84599984, -0.070495784, -1.3681931, 23.326256, -0.91202664, -0.064800754, 10.1774235, 22.84837, -0.9745514, -0.05906008, 21.472502, 22.32446, -1.033491, -0.053288586, 32.494568, 21.756693, -1.0887729, -0.04750085, 43.222256, 21.147306, -1.1403345, -0.041711222, 53.635315, 20.498589, -1.1881237, -0.035933767, 63.714672, 19.812881, -1.2320986, -0.030182252},
		'{220.94467, -22.134588, -0.68327236, 0.14565031, 209.72185, -22.745558, -0.58000046, 0.14303371, 198.2103, -23.28945, -0.4773432, 0.14012164, 186.44359, -23.766256, -0.3755374, 0.13692695, 174.4552, -24.176136, -0.27481315, 0.1334629, 162.27855, -24.519405, -0.17539336, 0.12974317, 149.94682, -24.796534, -0.0774935, 0.12578177, 137.49294, -25.008144, 0.018678905, 0.12159303, 124.94948, -25.155006, 0.11292458, 0.11719154, 112.34858, -25.23803, 0.20505281, 0.11259214, 99.72192, -25.258263, 0.29488173, 0.10780984, 87.100586, -25.216887, 0.3822386, 0.10285982, 74.51508, -25.115202, 0.4669601, 0.09775735, 61.9952, -24.954641, 0.54889244, 0.09251777, 49.570004, -24.73674, 0.62789166, 0.08715648, 37.267746, -24.463152, 0.70382357, 0.08168884, 25.115845, -24.135626, 0.77656424, 0.0761302, 13.140806, -23.756014, 0.84599984, 0.070495784, 1.3681931, -23.326256, 0.91202664, 0.064800754, -10.1774235, -22.84837, 0.9745514, 0.05906008, -21.472502, -22.32446, 1.033491, 0.053288586, -32.494568, -21.756693, 1.0887729, 0.04750085, -43.222256, -21.147306, 1.1403345, 0.041711222, -53.635315, -20.498589, 1.1881237, 0.035933767, -63.714672, -19.812881, 1.2320986, 0.030182252},
		'{672.33044, -39.69634, 3.066378, -0.18078938, 652.6359, -39.08045, 3.0294678, -0.18150762, 633.25134, -38.45651, 2.9914224, -0.18201949, 614.18054, -37.8255, 2.9523318, -0.18233427, 595.4269, -37.188354, 2.912282, -0.18246095, 576.99304, -36.545963, 2.8713567, -0.1824083, 558.8816, -35.89919, 2.8296363, -0.18218485, 541.0945, -35.24885, 2.7871976, -0.18179886, 523.63324, -34.595737, 2.744115, -0.18125838, 506.49905, -33.940594, 2.70046, -0.18057121, 489.69284, -33.284145, 2.6563008, -0.17974496, 473.215, -32.627075, 2.6117032, -0.17878693, 457.06573, -31.970037, 2.5667305, -0.17770432, 441.24484, -31.313652, 2.5214431, -0.17650399, 425.75186, -30.658514, 2.4758987, -0.17519264, 410.58603, -30.005186, 2.430153, -0.17377679, 395.74628, -29.354204, 2.3842585, -0.1722627, 381.23135, -28.706076, 2.3382664, -0.17065646, 367.03964, -28.061283, 2.2922244, -0.16896392, 353.16943, -27.420277, 2.246179, -0.1671908, 339.61868, -26.783493, 2.2001743, -0.16534257, 326.38516, -26.151333, 2.1542516, -0.16342454, 313.4665, -25.52418, 2.108451, -0.1614418, 300.86008, -24.902393, 2.0628097, -0.15939933, 288.56314, -24.286312, 2.0173643, -0.15730187},
		'{-672.33044, 39.69634, -3.066378, 0.18078938, -652.6359, 39.08045, -3.0294678, 0.18150762, -633.25134, 38.45651, -2.9914224, 0.18201949, -614.18054, 37.8255, -2.9523318, 0.18233427, -595.4269, 37.188354, -2.912282, 0.18246095, -576.99304, 36.545963, -2.8713567, 0.1824083, -558.8816, 35.89919, -2.8296363, 0.18218485, -541.0945, 35.24885, -2.7871976, 0.18179886, -523.63324, 34.595737, -2.744115, 0.18125838, -506.49905, 33.940594, -2.70046, 0.18057121, -489.69284, 33.284145, -2.6563008, 0.17974496, -473.215, 32.627075, -2.6117032, 0.17878693, -457.06573, 31.970037, -2.5667305, 0.17770432, -441.24484, 31.313652, -2.5214431, 0.17650399, -425.75186, 30.658514, -2.4758987, 0.17519264, -410.58603, 30.005186, -2.430153, 0.17377679, -395.74628, 29.354204, -2.3842585, 0.1722627, -381.23135, 28.706076, -2.3382664, 0.17065646, -367.03964, 28.061283, -2.2922244, 0.16896392, -353.16943, 27.420277, -2.246179, 0.1671908, -339.61868, 26.783493, -2.2001743, 0.16534257, -326.38516, 26.151333, -2.1542516, 0.16342454, -313.4665, 25.52418, -2.108451, 0.1614418, -300.86008, 24.902393, -2.0628097, 0.15939933, -288.56314, 24.286312, -2.0173643, 0.15730187}};
	localparam real Fbr[0:3][0:99] = '{
		'{183.25674, -17.803015, -1.9955642, -0.02115994, 191.84448, -16.545134, -2.006414, -0.027916582, 199.79929, -15.271762, -2.0121887, -0.034473382, 207.11423, -13.98629, -2.0129735, -0.040818363, 213.78412, -12.69207, -2.0088646, -0.046940286, 219.80539, -11.392408, -1.9999676, -0.05282868, 225.17615, -10.090563, -1.9863975, -0.058473844, 229.89612, -8.78973, -1.9682786, -0.06386685, 233.96657, -7.493044, -1.945744, -0.068999566, 237.39035, -6.2035656, -1.9189346, -0.073864646, 240.17183, -4.924279, -1.8879989, -0.07845553, 242.31682, -3.6580853, -1.8530928, -0.08276646, 243.83257, -2.4077973, -1.8143785, -0.086792454, 244.7277, -1.1761336, -1.7720243, -0.090529345, 245.01224, 0.03428483, -1.7262039, -0.093973726, 244.69739, 1.2209402, -1.6770965, -0.09712297, 243.79565, 2.3814216, -1.6248852, -0.09997521, 242.32071, 3.5134282, -1.5697573, -0.10252937, 240.28734, 4.614774, -1.5119035, -0.10478506, 237.71138, 5.683389, -1.4515173, -0.10674267, 234.60973, 6.7173247, -1.3887947, -0.10840329, 231.00014, 7.714753, -1.3239331, -0.109768696, 226.90134, 8.673971, -1.2571319, -0.110841356, 222.33281, 9.593401, -1.1885909, -0.111624405, 217.3148, 10.471594, -1.11851, -0.1121216},
		'{183.25674, -17.803015, -1.9955642, -0.02115994, 191.84448, -16.545134, -2.006414, -0.027916582, 199.79929, -15.271762, -2.0121887, -0.034473382, 207.11423, -13.98629, -2.0129735, -0.040818363, 213.78412, -12.69207, -2.0088646, -0.046940286, 219.80539, -11.392408, -1.9999676, -0.05282868, 225.17615, -10.090563, -1.9863975, -0.058473844, 229.89612, -8.78973, -1.9682786, -0.06386685, 233.96657, -7.493044, -1.945744, -0.068999566, 237.39035, -6.2035656, -1.9189346, -0.073864646, 240.17183, -4.924279, -1.8879989, -0.07845553, 242.31682, -3.6580853, -1.8530928, -0.08276646, 243.83257, -2.4077973, -1.8143785, -0.086792454, 244.7277, -1.1761336, -1.7720243, -0.090529345, 245.01224, 0.03428483, -1.7262039, -0.093973726, 244.69739, 1.2209402, -1.6770965, -0.09712297, 243.79565, 2.3814216, -1.6248852, -0.09997521, 242.32071, 3.5134282, -1.5697573, -0.10252937, 240.28734, 4.614774, -1.5119035, -0.10478506, 237.71138, 5.683389, -1.4515173, -0.10674267, 234.60973, 6.7173247, -1.3887947, -0.10840329, 231.00014, 7.714753, -1.3239331, -0.109768696, 226.90134, 8.673971, -1.2571319, -0.110841356, 222.33281, 9.593401, -1.1885909, -0.111624405, 217.3148, 10.471594, -1.11851, -0.1121216},
		'{182.00656, -17.691608, -1.9211302, -0.2637629, 190.55325, -16.50202, -1.8158827, -0.2539327, 198.51532, -15.352927, -1.7138801, -0.2443255, 205.9128, -14.243513, -1.615066, -0.23493986, 212.7653, -13.172956, -1.5193839, -0.22577423, 219.09207, -12.14044, -1.4267766, -0.21682692, 224.91194, -11.145147, -1.3371872, -0.20809613, 230.24329, -10.186268, -1.2505579, -0.19957995, 235.10413, -9.262992, -1.1668315, -0.19127631, 239.51207, -8.374516, -1.0859503, -0.18318307, 243.48431, -7.520039, -1.0078568, -0.17529799, 247.03764, -6.6987696, -0.93249375, -0.16761872, 250.18848, -5.909919, -0.85980356, -0.16014284, 252.95282, -5.1527047, -0.7897292, -0.15286785, 255.34631, -4.4263535, -0.7222136, -0.14579117, 257.3842, -3.7300978, -0.6572003, -0.13891017, 259.0813, -3.0631773, -0.5946326, -0.13222215, 260.45212, -2.4248407, -0.5344547, -0.12572433, 261.51077, -1.8143445, -0.47661078, -0.11941391, 262.27097, -1.2309542, -0.42104563, -0.11328804, 262.74612, -0.67394376, -0.36770442, -0.10734382, 262.9492, -0.14259684, -0.3165328, -0.10157833, 262.89285, 0.3637938, -0.26747695, -0.095988594, 262.58945, 0.84592545, -0.22048353, -0.09057163, 262.05087, 1.3044858, -0.17549983, -0.08532442},
		'{182.00656, -17.691608, -1.9211302, -0.2637629, 190.55325, -16.50202, -1.8158827, -0.2539327, 198.51532, -15.352927, -1.7138801, -0.2443255, 205.9128, -14.243513, -1.615066, -0.23493986, 212.7653, -13.172956, -1.5193839, -0.22577423, 219.09207, -12.14044, -1.4267766, -0.21682692, 224.91194, -11.145147, -1.3371872, -0.20809613, 230.24329, -10.186268, -1.2505579, -0.19957995, 235.10413, -9.262992, -1.1668315, -0.19127631, 239.51207, -8.374516, -1.0859503, -0.18318307, 243.48431, -7.520039, -1.0078568, -0.17529799, 247.03764, -6.6987696, -0.93249375, -0.16761872, 250.18848, -5.909919, -0.85980356, -0.16014284, 252.95282, -5.1527047, -0.7897292, -0.15286785, 255.34631, -4.4263535, -0.7222136, -0.14579117, 257.3842, -3.7300978, -0.6572003, -0.13891017, 259.0813, -3.0631773, -0.5946326, -0.13222215, 260.45212, -2.4248407, -0.5344547, -0.12572433, 261.51077, -1.8143445, -0.47661078, -0.11941391, 262.27097, -1.2309542, -0.42104563, -0.11328804, 262.74612, -0.67394376, -0.36770442, -0.10734382, 262.9492, -0.14259684, -0.3165328, -0.10157833, 262.89285, 0.3637938, -0.26747695, -0.095988594, 262.58945, 0.84592545, -0.22048353, -0.09057163, 262.05087, 1.3044858, -0.17549983, -0.08532442}};
	localparam real Fbi[0:3][0:99] = '{
		'{-220.94467, -22.134588, 0.68327236, 0.14565031, -209.72185, -22.745558, 0.58000046, 0.14303371, -198.2103, -23.28945, 0.4773432, 0.14012164, -186.44359, -23.766256, 0.3755374, 0.13692695, -174.4552, -24.176136, 0.27481315, 0.1334629, -162.27855, -24.519405, 0.17539336, 0.12974317, -149.94682, -24.796534, 0.0774935, 0.12578177, -137.49294, -25.008144, -0.018678905, 0.12159303, -124.94948, -25.155006, -0.11292458, 0.11719154, -112.34858, -25.23803, -0.20505281, 0.11259214, -99.72192, -25.258263, -0.29488173, 0.10780984, -87.100586, -25.216887, -0.3822386, 0.10285982, -74.51508, -25.115202, -0.4669601, 0.09775735, -61.9952, -24.954641, -0.54889244, 0.09251777, -49.570004, -24.73674, -0.62789166, 0.08715648, -37.267746, -24.463152, -0.70382357, 0.08168884, -25.115845, -24.135626, -0.77656424, 0.0761302, -13.140806, -23.756014, -0.84599984, 0.070495784, -1.3681931, -23.326256, -0.91202664, 0.064800754, 10.1774235, -22.84837, -0.9745514, 0.05906008, 21.472502, -22.32446, -1.033491, 0.053288586, 32.494568, -21.756693, -1.0887729, 0.04750085, 43.222256, -21.147306, -1.1403345, 0.041711222, 53.635315, -20.498589, -1.1881237, 0.035933767, 63.714672, -19.812881, -1.2320986, 0.030182252},
		'{220.94467, 22.134588, -0.68327236, -0.14565031, 209.72185, 22.745558, -0.58000046, -0.14303371, 198.2103, 23.28945, -0.4773432, -0.14012164, 186.44359, 23.766256, -0.3755374, -0.13692695, 174.4552, 24.176136, -0.27481315, -0.1334629, 162.27855, 24.519405, -0.17539336, -0.12974317, 149.94682, 24.796534, -0.0774935, -0.12578177, 137.49294, 25.008144, 0.018678905, -0.12159303, 124.94948, 25.155006, 0.11292458, -0.11719154, 112.34858, 25.23803, 0.20505281, -0.11259214, 99.72192, 25.258263, 0.29488173, -0.10780984, 87.100586, 25.216887, 0.3822386, -0.10285982, 74.51508, 25.115202, 0.4669601, -0.09775735, 61.9952, 24.954641, 0.54889244, -0.09251777, 49.570004, 24.73674, 0.62789166, -0.08715648, 37.267746, 24.463152, 0.70382357, -0.08168884, 25.115845, 24.135626, 0.77656424, -0.0761302, 13.140806, 23.756014, 0.84599984, -0.070495784, 1.3681931, 23.326256, 0.91202664, -0.064800754, -10.1774235, 22.84837, 0.9745514, -0.05906008, -21.472502, 22.32446, 1.033491, -0.053288586, -32.494568, 21.756693, 1.0887729, -0.04750085, -43.222256, 21.147306, 1.1403345, -0.041711222, -53.635315, 20.498589, 1.1881237, -0.035933767, -63.714672, 19.812881, 1.2320986, -0.030182252},
		'{-672.33044, -39.69634, -3.066378, -0.18078938, -652.6359, -39.08045, -3.0294678, -0.18150762, -633.25134, -38.45651, -2.9914224, -0.18201949, -614.18054, -37.8255, -2.9523318, -0.18233427, -595.4269, -37.188354, -2.912282, -0.18246095, -576.99304, -36.545963, -2.8713567, -0.1824083, -558.8816, -35.89919, -2.8296363, -0.18218485, -541.0945, -35.24885, -2.7871976, -0.18179886, -523.63324, -34.595737, -2.744115, -0.18125838, -506.49905, -33.940594, -2.70046, -0.18057121, -489.69284, -33.284145, -2.6563008, -0.17974496, -473.215, -32.627075, -2.6117032, -0.17878693, -457.06573, -31.970037, -2.5667305, -0.17770432, -441.24484, -31.313652, -2.5214431, -0.17650399, -425.75186, -30.658514, -2.4758987, -0.17519264, -410.58603, -30.005186, -2.430153, -0.17377679, -395.74628, -29.354204, -2.3842585, -0.1722627, -381.23135, -28.706076, -2.3382664, -0.17065646, -367.03964, -28.061283, -2.2922244, -0.16896392, -353.16943, -27.420277, -2.246179, -0.1671908, -339.61868, -26.783493, -2.2001743, -0.16534257, -326.38516, -26.151333, -2.1542516, -0.16342454, -313.4665, -25.52418, -2.108451, -0.1614418, -300.86008, -24.902393, -2.0628097, -0.15939933, -288.56314, -24.286312, -2.0173643, -0.15730187},
		'{672.33044, 39.69634, 3.066378, 0.18078938, 652.6359, 39.08045, 3.0294678, 0.18150762, 633.25134, 38.45651, 2.9914224, 0.18201949, 614.18054, 37.8255, 2.9523318, 0.18233427, 595.4269, 37.188354, 2.912282, 0.18246095, 576.99304, 36.545963, 2.8713567, 0.1824083, 558.8816, 35.89919, 2.8296363, 0.18218485, 541.0945, 35.24885, 2.7871976, 0.18179886, 523.63324, 34.595737, 2.744115, 0.18125838, 506.49905, 33.940594, 2.70046, 0.18057121, 489.69284, 33.284145, 2.6563008, 0.17974496, 473.215, 32.627075, 2.6117032, 0.17878693, 457.06573, 31.970037, 2.5667305, 0.17770432, 441.24484, 31.313652, 2.5214431, 0.17650399, 425.75186, 30.658514, 2.4758987, 0.17519264, 410.58603, 30.005186, 2.430153, 0.17377679, 395.74628, 29.354204, 2.3842585, 0.1722627, 381.23135, 28.706076, 2.3382664, 0.17065646, 367.03964, 28.061283, 2.2922244, 0.16896392, 353.16943, 27.420277, 2.246179, 0.1671908, 339.61868, 26.783493, 2.2001743, 0.16534257, 326.38516, 26.151333, 2.1542516, 0.16342454, 313.4665, 25.52418, 2.108451, 0.1614418, 300.86008, 24.902393, 2.0628097, 0.15939933, 288.56314, 24.286312, 2.0173643, 0.15730187}};
	localparam real hf[0:1199] = {0.016714763, -1.6967899e-05, -2.2033028e-05, 4.3969756e-08, 0.016697802, -5.0869214e-05, -2.1941874e-05, 1.316649e-07, 0.01666391, -8.466729e-05, -2.1759943e-05, 2.1863927e-07, 0.016613163, -0.00011829375, -2.148794e-05, 3.0443857e-07, 0.016545657, -0.00015168074, -2.1126889e-05, 3.886314e-07, 0.016461533, -0.00018476119, -2.0678113e-05, 4.7080962e-07, 0.016360957, -0.00021746896, -2.0143225e-05, 5.505885e-07, 0.016244136, -0.00024973904, -1.9524112e-05, 6.276069e-07, 0.016111301, -0.00028150773, -1.8822926e-05, 7.0152754e-07, 0.015962722, -0.00031271283, -1.8042067e-05, 7.7203686e-07, 0.015798694, -0.00034329374, -1.7184168e-05, 8.3884527e-07, 0.0156195415, -0.00037319172, -1.6252085e-05, 9.016869e-07, 0.015425624, -0.00040234992, -1.5248873e-05, 9.603198e-07, 0.015217324, -0.00043071364, -1.41777855e-05, 1.0145253e-06, 0.014995052, -0.00045823032, -1.3042247e-05, 1.0641085e-06, 0.0147592435, -0.0004848498, -1.1845846e-05, 1.1088973e-06, 0.01451036, -0.0005105243, -1.0592313e-05, 1.1487429e-06, 0.014248883, -0.0005352087, -9.285516e-06, 1.1835186e-06, 0.013975322, -0.0005588603, -7.929435e-06, 1.2131203e-06, 0.013690202, -0.0005814394, -6.5281547e-06, 1.2374652e-06, 0.013394068, -0.00060290896, -5.0858453e-06, 1.2564922e-06, 0.013087483, -0.0006232347, -3.6067513e-06, 1.2701607e-06, 0.012771029, -0.00064238557, -2.0951757e-06, 1.2784507e-06, 0.012445298, -0.0006603331, -5.554659e-07, 1.2813616e-06, 0.0121109, -0.0006770521, 1.0079999e-06, 1.278912e-06, 0.011768455, -0.00069252035, 2.590826e-06, 1.271139e-06, 0.011418591, -0.00070671865, 4.188613e-06, 1.2580974e-06, 0.011061951, -0.0007196309, 5.7969696e-06, 1.2398594e-06, 0.010699177, -0.00073124404, 7.4115273e-06, 1.2165135e-06, 0.010330924, -0.00074154814, 9.02795e-06, 1.1881637e-06, 0.009957848, -0.0007505362, 1.0641949e-05, 1.154929e-06, 0.0095806075, -0.00075820443, 1.2249292e-05, 1.1169429e-06, 0.009199864, -0.0007645519, 1.3845814e-05, 1.0743521e-06, 0.008816276, -0.0007695808, 1.5427428e-05, 1.0273158e-06, 0.008430502, -0.00077329593, 1.699014e-05, 9.760051e-07, 0.008043197, -0.0007757053, 1.8530049e-05, 9.2060213e-07, 0.0076550124, -0.0007768197, 2.0043366e-05, 8.612991e-07, 0.0072665913, -0.0007766524, 2.1526417e-05, 7.982977e-07, 0.006878571, -0.0007752197, 2.2975652e-05, 7.318081e-07, 0.0064915796, -0.0007725403, 2.4387655e-05, 6.6204797e-07, 0.006106235, -0.0007686354, 2.5759146e-05, 5.892422e-07, 0.0057231444, -0.00076352886, 2.7086993e-05, 5.1362133e-07, 0.005342902, -0.0007572467, 2.8368218e-05, 4.3542153e-07, 0.004966089, -0.0007498172, 2.96e-05, 3.5488307e-07, 0.004593271, -0.00074127084, 3.0779676e-05, 2.7225e-07, 0.004224999, -0.0007316402, 3.1904754e-05, 1.8776915e-07, 0.003861806, -0.0007209598, 3.2972916e-05, 1.016894e-07, 0.003504208, -0.00070926594, 3.3982007e-05, 1.4260949e-08, 0.0031527025, -0.00069659663, 3.4930064e-05, -7.4265515e-08, 0.0028077674, -0.0006829916, 3.5815297e-05, -1.6363948e-07, 0.00246986, -0.0006684919, 3.663609e-05, -2.5361132e-07, 0.0021394175, -0.0006531401, 3.7391026e-05, -3.4393307e-07, 0.0018168548, -0.00063697994, 3.8078855e-05, -4.3435898e-07, 0.0015025649, -0.0006200564, 3.869852e-05, -5.246463e-07, 0.0011969181, -0.00060241536, 3.9249146e-05, -6.145557e-07, 0.0009002614, -0.0005841035, 3.973004e-05, -7.0385215e-07, 0.00061291846, -0.0005651685, 4.0140687e-05, -7.9230534e-07, 0.0003351888, -0.0005456585, 4.048076e-05, -8.796902e-07, 6.734773e-05, -0.0005256222, 4.0750107e-05, -9.657875e-07, -0.00019035382, -0.00050510874, 4.0948744e-05, -1.0503844e-06, -0.00043768962, -0.0004841674, 4.1076873e-05, -1.1332747e-06, -0.0006744581, -0.00046284776, 4.113486e-05, -1.2142597e-06, -0.0009004825, -0.00044119937, 4.112323e-05, -1.293148e-06, -0.0011156108, -0.00041927173, 4.1042673e-05, -1.3697564e-06, -0.0013197159, -0.00039711408, 4.0894043e-05, -1.4439103e-06, -0.0015126948, -0.0003747754, 4.0678347e-05, -1.5154434e-06, -0.0016944691, -0.00035230428, 4.0396728e-05, -1.5841987e-06, -0.0018649849, -0.00032974873, 4.005048e-05, -1.6500285e-06, -0.0020242117, -0.0003071562, 3.9641036e-05, -1.7127944e-06, -0.0021721425, -0.00028457335, 3.9169958e-05, -1.7723679e-06, -0.0023087943, -0.00026204612, 3.8638926e-05, -1.8286304e-06, -0.0024342055, -0.00023961939, 3.804975e-05, -1.8814732e-06, -0.0025484376, -0.00021733719, 3.7404352e-05, -1.9307977e-06, -0.0026515739, -0.00019524238, 3.670475e-05, -1.976516e-06, -0.0027437182, -0.00017337665, 3.5953068e-05, -2.0185496e-06, -0.0028249954, -0.00015178052, 3.5151523e-05, -2.0568316e-06, -0.00289555, -0.00013049312, 3.430242e-05, -2.0913042e-06, -0.0029555461, -0.000109552224, 3.3408134e-05, -2.1219207e-06, -0.003005166, -8.899417e-05, 3.2471118e-05, -2.1486442e-06, -0.00304461, -6.8853784e-05, 3.149389e-05, -2.1714486e-06, -0.003074095, -4.9164333e-05, 3.0479021e-05, -2.1903172e-06, -0.0030938545, -2.9957473e-05, 2.9429133e-05, -2.2052434e-06, -0.0031041377, -1.1263215e-05, 2.834689e-05, -2.216231e-06, -0.003105208, 6.8901313e-06, 2.7234997e-05, -2.2232928e-06, -0.0030973423, 2.447598e-05, 2.6096179e-05, -2.226451e-06, -0.0030808307, 4.1469506e-05, 2.4933186e-05, -2.2257375e-06, -0.0030559753, 5.7847665e-05, 2.3748784e-05, -2.2211932e-06, -0.0030230891, 7.3589224e-05, 2.2545744e-05, -2.2128672e-06, -0.0029824954, 8.8674766e-05, 2.1326836e-05, -2.2008176e-06, -0.0029345267, 0.00010308671, 2.0094829e-05, -2.1851106e-06, -0.0028795234, 0.00011680934, 1.8852472e-05, -2.16582e-06, -0.0028178345, 0.00012982874, 1.7602502e-05, -2.1430276e-06, -0.002749814, 0.00014213285, 1.6347625e-05, -2.1168223e-06, -0.0026758225, 0.00015371149, 1.5090519e-05, -2.0872997e-06, -0.002596225, 0.00016455624, 1.3833823e-05, -2.0545624e-06, -0.0025113896, 0.00017466056, 1.2580132e-05, -2.0187185e-06, -0.0024216885, 0.00018401962, 1.1331994e-05, -1.9798829e-06, -0.0023274948, 0.00019263044, 1.0091903e-05, -1.938175e-06, -0.002229183, 0.00020049176, 8.8622955e-06, -1.8937199e-06, -0.002127128, 0.00020760401, 7.64554e-06, -1.846647e-06, -0.0020217034, 0.00021396932, 6.443941e-06, -1.7970901e-06, -0.0019132824, 0.0002195915, 5.2597284e-06, -1.745187e-06, -0.0018022349, 0.0002244759, 4.0950563e-06, -1.6910788e-06, -0.0016889283, 0.00022862946, 2.9519979e-06, -1.6349095e-06, -0.001573726, 0.00023206066, 1.8325427e-06, -1.5768263e-06, -0.0014569864, 0.00023477942, 7.38593e-07, -1.5169782e-06, -0.0013390634, 0.0002367971, -3.2803908e-07, -1.4555162e-06, -0.001220304, 0.00023812639, -1.3656344e-06, -1.3925928e-06, -0.0011010494, 0.00023878133, -2.372569e-06, -1.3283615e-06, -0.0009816326, 0.00023877717, -3.3473168e-06, -1.2629763e-06, -0.0008623794, 0.00023813036, -4.288451e-06, -1.1965919e-06, -0.0007436065, 0.0002368585, -5.1946454e-06, -1.1293628e-06, -0.000625622, 0.00023498024, -6.0646767e-06, -1.0614427e-06, -0.0005087241, 0.00023251523, -6.897425e-06, -9.929848e-07, -0.00039320113, 0.00022948405, -7.691875e-06, -9.24141e-07, -0.00027933085, 0.00022590818, -8.447116e-06, -8.550617e-07, -0.00016738006, 0.00022180987, -9.162341e-06, -7.858955e-07, -5.7604266e-05, 0.0002172121, -9.83685e-06, -7.1678863e-07, 4.9752703e-05, 0.00021213855, -1.0470048e-05, -6.4788503e-07, 0.00015445899, 0.00020661348, -1.1061443e-05, -5.7932573e-07, 0.00025629502, 0.00020066166, -1.1610647e-05, -5.1124863e-07, 0.0003550537, 0.00019430835, -1.2117375e-05, -4.437883e-07, 0.00045054068, 0.0001875792, -1.2581445e-05, -3.7707576e-07, 0.00054257456, 0.00018050017, -1.3002771e-05, -3.11238e-07, 0.0006309869, 0.00017309746, -1.338137e-05, -2.46398e-07, 0.00071562245, 0.00016539752, -1.3717353e-05, -1.826743e-07, 0.00079633924, 0.00015742687, -1.4010926e-05, -1.2018099e-07, 0.00087300857, 0.0001492121, -1.4262389e-05, -5.9027336e-08, 0.00094551506, 0.0001407798, -1.447213e-05, 6.822579e-10, 0.0010137565, 0.0001321565, -1.4640624e-05, 5.8848492e-08, 0.0010776441, 0.00012336859, -1.4768433e-05, 1.153773e-07, 0.001137102, 0.00011444229, -1.4856199e-05, 1.7017996e-07, 0.0011920676, 0.000105403546, -1.4904645e-05, 2.2317325e-07, 0.0012424911, 9.627802e-05, -1.4914564e-05, 2.7427947e-07, 0.0012883353, 8.7091015e-05, -1.4886829e-05, 3.2342666e-07, 0.0013295759, 7.7867415e-05, -1.4822377e-05, 3.7054852e-07, 0.0013662007, 6.863166e-05, -1.4722211e-05, 4.1558457e-07, 0.0013982096, 5.940767e-05, -1.4587396e-05, 4.5848014e-07, 0.0014256142, 5.0218805e-05, -1.4419057e-05, 4.991864e-07, 0.001448438, 4.108784e-05, -1.4218371e-05, 5.3766047e-07, 0.0014667154, 3.203689e-05, -1.3986567e-05, 5.7386524e-07, 0.0014804917, 2.3087405e-05, -1.3724919e-05, 6.077694e-07, 0.0014898231, 1.4260112e-05, -1.34347465e-05, 6.3934755e-07, 0.0014947755, 5.5749824e-06, -1.3117407e-05, 6.6857996e-07, 0.001495425, -2.948796e-06, -1.27742915e-05, 6.9545274e-07, 0.0014918568, -1.1292848e-05, -1.2406825e-05, 7.199574e-07, 0.001484165, -1.9439643e-05, -1.2016456e-05, 7.4209134e-07, 0.0014724527, -2.7372516e-05, -1.1604659e-05, 7.6185705e-07, 0.0014568308, -3.507569e-05, -1.1172928e-05, 7.7926256e-07, 0.0014374178, -4.253429e-05, -1.072277e-05, 7.943212e-07, 0.0014143395, -4.973438e-05, -1.0255704e-05, 8.070512e-07, 0.0013877286, -5.666295e-05, -9.77326e-06, 8.1747595e-07, 0.0013577238, -6.330795e-05, -9.276969e-06, 8.2562354e-07, 0.0013244698, -6.965827e-05, -8.768362e-06, 8.3152685e-07, 0.0012881164, -7.570381e-05, -8.248969e-06, 8.3522303e-07, 0.0012488184, -8.143539e-05, -7.72031e-06, 8.3675377e-07, 0.0012067347, -8.684485e-05, -7.1838986e-06, 8.361648e-07, 0.0011620284, -9.1924965e-05, -6.641231e-06, 8.33506e-07, 0.0011148656, -9.66695e-05, -6.093788e-06, 8.288307e-07, 0.0010654157, -0.000101073194, -5.543032e-06, 8.221961e-07, 0.00101385, -0.000105131716, -4.9903992e-06, 8.1366267e-07, 0.00096034206, -0.00010884172, -4.4373014e-06, 8.032939e-07, 0.0009050668, -0.00011220076, -3.8851213e-06, 7.9115654e-07, 0.00084820006, -0.000115207346, -3.3352094e-06, 7.7731977e-07, 0.0007899183, -0.00011786087, -2.7888827e-06, 7.618556e-07, 0.000730398, -0.00012016164, -2.2474212e-06, 7.448381e-07, 0.0006698153, -0.00012211081, -1.7120661e-06, 7.263435e-07, 0.0006083455, -0.00012371042, -1.1840173e-06, 7.0645007e-07, 0.0005461627, -0.0001249633, -6.6443147e-07, 6.8523747e-07, 0.0004834394, -0.0001258731, -1.544205e-07, 6.6278704e-07, 0.00042034604, -0.00012644428, 3.4495065e-07, 6.391811e-07, 0.0003570507, -0.000126682, 8.3266536e-07, 6.145032e-07, 0.00029371865, -0.00012659217, 1.3077569e-06, 5.888375e-07, 0.00023051204, -0.0001261814, 1.7693094e-06, 5.622688e-07, 0.00016758955, -0.00012545697, 2.2164597e-06, 5.348822e-07, 0.00010510606, -0.00012442676, 2.6483974e-06, 5.0676306e-07, 4.3212363e-05, -0.00012309928, 3.0643669e-06, 4.7799654e-07, -1.7945164e-05, -0.000121483616, 3.4636669e-06, 4.4866758e-07, -7.8224795e-05, -0.00011958936, 3.8456515e-06, 4.188608e-07, -0.00013748975, -0.00011742662, 4.2097313e-06, 3.8866e-07, -0.0001956084, -0.00011500597, 4.555372e-06, 3.5814827e-07, -0.00025245454, -0.0001123384, 4.8820966e-06, 3.274076e-07, -0.00030790752, -0.000109435314, 5.189484e-06, 2.9651886e-07, -0.00036185252, -0.000106308464, 5.4771685e-06, 2.6556154e-07, -0.0004141807, -0.00010296991, 5.7448415e-06, 2.3461364e-07, -0.0004647892, -9.943203e-05, 5.9922486e-06, 2.0375144e-07, -0.00051358156, -9.5707415e-05, 6.219192e-06, 1.7304944e-07, -0.0005604676, -9.1808906e-05, 6.425527e-06, 1.425802e-07, -0.00060536363, -8.774949e-05, 6.611162e-06, 1.1241415e-07, -0.0006481924, -8.354231e-05, 6.7760593e-06, 8.2619515e-08, -0.0006888835, -7.9200625e-05, 6.9202333e-06, 5.326218e-08, -0.0007273728, -7.473775e-05, 7.043747e-06, 2.4405603e-08, -0.00076360325, -7.016705e-05, 7.1467143e-06, -3.889324e-09, -0.0007975241, -6.5501896e-05, 7.2292974e-06, -3.1564344e-08, -0.0008290916, -6.075562e-05, 7.291704e-06, -5.856393e-08, -0.0008582684, -5.5941502e-05, 7.3341894e-06, -8.483536e-08, -0.00088502397, -5.107273e-05, 7.3570504e-06, -1.1032878e-07, -0.0009093342, -4.616237e-05, 7.3606266e-06, -1.3499728e-07, -0.00093118154, -4.1223335e-05, 7.3452993e-06, -1.5879695e-07, -0.00095055485, -3.6268357e-05, 7.311487e-06, -1.8168689e-07, -0.00096744933, -3.130996e-05, 7.2596463e-06, -2.0362927e-07, -0.0009818663, -2.6360438e-05, 7.1902678e-06, -2.245894e-07, -0.0009938133, -2.1431819e-05, 7.1038767e-06, -2.4453567e-07, -0.0010033036, -1.653585e-05, 7.001028e-06, -2.634396e-07, -0.0010103564, -1.1683969e-05, 6.882307e-06, -2.8127587e-07, -0.0010149967, -6.887285e-06, 6.7483256e-06, -2.9802231e-07, -0.0010172547, -2.1565565e-06, 6.5997215e-06, -3.1365983e-07, -0.001017166, 2.4978276e-06, 6.437155e-06, -3.2817246e-07, -0.0010147712, 7.0658666e-06, 6.261308e-06, -3.4154735e-07, -0.0010101161, 1.1537964e-05, 6.0728808e-06, -3.5377462e-07, -0.0010032507, 1.5904945e-05, 5.872591e-06, -3.6484752e-07, -0.00099423, 2.0158068e-05, 5.6611707e-06, -3.7476218e-07, -0.0009831131, 2.4289038e-05, 5.4393654e-06, -3.8351766e-07, -0.0009699627, 2.8290024e-05, 5.2079304e-06, -3.9111592e-07, -0.0009548459, 3.2153654e-05, 4.9676296e-06, -3.9756165e-07, -0.0009378331, 3.5873047e-05, 4.7192348e-06, -4.0286236e-07, -0.000918998, 3.94418e-05, 4.463521e-06, -4.0702812e-07, -0.0008984174, 4.2853997e-05, 4.2012653e-06, -4.1007166e-07, -0.00087617093, 4.610423e-05, 3.933247e-06, -4.1200818e-07, -0.00085234095, 4.918758e-05, 3.660244e-06, -4.1285523e-07, -0.00082701194, 5.2099636e-05, 3.383029e-06, -4.1263277e-07, -0.0008002705, 5.4836495e-05, 3.1023721e-06, -4.113629e-07, -0.0007722052, 5.7394747e-05, 2.8190354e-06, -4.090699e-07, -0.000742906, 5.9771486e-05, 2.5337724e-06, -4.0578007e-07, -0.0007124644, 6.196431e-05, 2.2473273e-06, -4.015216e-07, -0.0006809727, 6.397131e-05, 1.9604315e-06, -3.9632445e-07, -0.00064852426, 6.5791064e-05, 1.6738037e-06, -3.9022038e-07, -0.000615213, 6.742264e-05, 1.3881476e-06, -3.8324262e-07, -0.00058113306, 6.8865564e-05, 1.1041507e-06, -3.7542603e-07, -0.0005463789, 7.011986e-05, 8.224829e-07, -3.6680666e-07, -0.0005110446, 7.118599e-05, 5.437951e-07, -3.574219e-07, -0.0004752241, 7.206488e-05, 2.6871828e-07, -3.4731028e-07, -0.0004390107, 7.275787e-05, -2.1380147e-09, -3.365113e-07, -0.00040249692, 7.326677e-05, -2.6818645e-07, -3.250654e-07, -0.00036577426, 7.359374e-05, -5.2886304e-07, -3.1301374e-07, -0.00032893306, 7.3741416e-05, -7.8362797e-07, -3.003982e-07, -0.00029206224, 7.3712756e-05, -1.0319665e-06, -2.8726117e-07, -0.00025524915, 7.351113e-05, -1.2733898e-06, -2.7364553e-07, -0.00021857933, 7.314025e-05, -1.5074353e-06, -2.5959437e-07, -0.00018213644, 7.2604154e-05, -1.7336679e-06, -2.4515114e-07, -0.000146002, 7.1907234e-05, -1.95168e-06, -2.303593e-07, -0.00011025524, 7.105417e-05, -2.1610917e-06, -2.1526229e-07, -7.497303e-05, 7.004994e-05, -2.361552e-06, -1.9990347e-07, -4.022964e-05, 6.889978e-05, -2.552739e-06, -1.8432597e-07, -6.096666e-06, 6.7609195e-05, -2.7343588e-06, -1.6857263e-07, 2.7357097e-05, 6.618392e-05, -2.9061473e-06, -1.5268581e-07, 6.0065784e-05, 6.462991e-05, -3.0678696e-06, -1.3670744e-07, 9.196656e-05, 6.295331e-05, -3.2193198e-06, -1.2067878e-07, 0.0001229997, 6.116045e-05, -3.360321e-06, -1.0464043e-07, 0.0001531087, 5.925783e-05, -3.4907257e-06, -8.86322e-08, 0.00018224033, 5.7252073e-05, -3.6104145e-06, -7.2693055e-08, 0.0002103447, 5.514994e-05, -3.7192976e-06, -5.686101e-08, 0.00023737534, 5.295829e-05, -3.817312e-06, -4.1173067e-08, 0.00026328923, 5.0684073e-05, -3.904424e-06, -2.5665162e-08, 0.0002880468, 4.8334296e-05, -3.9806255e-06, -1.037207e-08, 0.0003116121, 4.591602e-05, -4.0459363e-06, 4.67264e-09, 0.00033395257, 4.343634e-05, -4.1004023e-06, 1.9436667e-08, 0.00035503937, 4.090236e-05, -4.1440944e-06, 3.388903e-08, 0.00037484706, 3.832118e-05, -4.1771095e-06, 4.800012e-08, 0.00039335384, 3.5699883e-05, -4.1995677e-06, 6.1741744e-08, 0.00041054143, 3.30455e-05, -4.211613e-06, 7.508717e-08, 0.00042639498, 3.0365021e-05, -4.213412e-06, 8.801115e-08, 0.00044090324, 2.7665357e-05, -4.2051524e-06, 1.0048996e-07, 0.0004540583, 2.4953339e-05, -4.187044e-06, 1.1250146e-07, 0.0004658556, 2.2235692e-05, -4.1593153e-06, 1.2402504e-07, 0.00047629414, 1.9519026e-05, -4.1222147e-06, 1.350417e-07, 0.0004853759, 1.6809823e-05, -4.0760087e-06, 1.4553409e-07, 0.00049310626, 1.4114422e-05, -4.02098e-06, 1.5548643e-07, 0.0004994936, 1.1439008e-05, -3.9574284e-06, 1.648846e-07, 0.0005045496, 8.789597e-06, -3.8856674e-06, 1.7371607e-07, 0.0005082885, 6.172028e-06, -3.8060255e-06, 1.8197001e-07, 0.00051072787, 3.5919504e-06, -3.7188438e-06, 1.8963712e-07, 0.00051188766, 1.054814e-06, -3.624475e-06, 1.9670982e-07, 0.0005117907, -1.4341393e-06, -3.5232827e-06, 2.0318203e-07, 0.0005104623, -3.8698854e-06, -3.4156399e-06, 2.0904932e-07, 0.00050793047, -6.2476247e-06, -3.3019278e-06, 2.143088e-07, 0.00050422514, -8.562791e-06, -3.182536e-06, 2.1895912e-07, 0.00049937883, -1.0811055e-05, -3.0578592e-06, 2.2300044e-07, 0.00049342593, -1.2988336e-05, -2.928298e-06, 2.2643444e-07, 0.00048640295, -1.5090798e-05, -2.7942576e-06, 2.2926419e-07, 0.0004783482, -1.7114864e-05, -2.6561452e-06, 2.3149421e-07, 0.0004693017, -1.9057215e-05, -2.5143706e-06, 2.331304e-07, 0.0004593051, -2.091479e-05, -2.369345e-06, 2.3417998e-07, 0.0004484015, -2.2684793e-05, -2.221479e-06, 2.3465147e-07, 0.00043663534, -2.4364694e-05, -2.0711823e-06, 2.3455462e-07, 0.0004240522, -2.5952228e-05, -1.9188628e-06, 2.3390038e-07, 0.00041069882, -2.7445398e-05, -1.7649253e-06, 2.3270088e-07, 0.0003966228, -2.8842473e-05, -1.6097708e-06, 2.309693e-07, 0.0003818726, -3.0141984e-05, -1.4537956e-06, 2.2871988e-07, 0.0003664973, -3.134273e-05, -1.2973902e-06, 2.2596784e-07, 0.0003505465, -3.244377e-05, -1.1409387e-06, 2.2272935e-07, 0.00033407027, -3.344442e-05, -9.84818e-07, 2.1902143e-07, 0.0003171189, -3.434425e-05, -8.293968e-07, 2.1486191e-07, 0.00029974285, -3.514309e-05, -6.750352e-07, 2.102694e-07, 0.00028199263, -3.5841003e-05, -5.2208367e-07, 2.0526318e-07, 0.00026391863, -3.6438305e-05, -3.7088242e-07, 1.998632e-07, 0.000245571, -3.6935544e-05, -2.2176111e-07, 1.940899e-07, 0.00022699962, -3.7333502e-05, -7.5037846e-08, 1.8796436e-07, 0.00020825388, -3.7633177e-05, 6.8981144e-08, 1.81508e-07, 0.00018938263, -3.7835795e-05, 2.1000207e-07, 1.7474268e-07};
	localparam real hb[0:1199] = {0.016714763, 1.6967899e-05, -2.2033028e-05, -4.3969756e-08, 0.016697802, 5.0869214e-05, -2.1941874e-05, -1.316649e-07, 0.01666391, 8.466729e-05, -2.1759943e-05, -2.1863927e-07, 0.016613163, 0.00011829375, -2.148794e-05, -3.0443857e-07, 0.016545657, 0.00015168074, -2.1126889e-05, -3.886314e-07, 0.016461533, 0.00018476119, -2.0678113e-05, -4.7080962e-07, 0.016360957, 0.00021746896, -2.0143225e-05, -5.505885e-07, 0.016244136, 0.00024973904, -1.9524112e-05, -6.276069e-07, 0.016111301, 0.00028150773, -1.8822926e-05, -7.0152754e-07, 0.015962722, 0.00031271283, -1.8042067e-05, -7.7203686e-07, 0.015798694, 0.00034329374, -1.7184168e-05, -8.3884527e-07, 0.0156195415, 0.00037319172, -1.6252085e-05, -9.016869e-07, 0.015425624, 0.00040234992, -1.5248873e-05, -9.603198e-07, 0.015217324, 0.00043071364, -1.41777855e-05, -1.0145253e-06, 0.014995052, 0.00045823032, -1.3042247e-05, -1.0641085e-06, 0.0147592435, 0.0004848498, -1.1845846e-05, -1.1088973e-06, 0.01451036, 0.0005105243, -1.0592313e-05, -1.1487429e-06, 0.014248883, 0.0005352087, -9.285516e-06, -1.1835186e-06, 0.013975322, 0.0005588603, -7.929435e-06, -1.2131203e-06, 0.013690202, 0.0005814394, -6.5281547e-06, -1.2374652e-06, 0.013394068, 0.00060290896, -5.0858453e-06, -1.2564922e-06, 0.013087483, 0.0006232347, -3.6067513e-06, -1.2701607e-06, 0.012771029, 0.00064238557, -2.0951757e-06, -1.2784507e-06, 0.012445298, 0.0006603331, -5.554659e-07, -1.2813616e-06, 0.0121109, 0.0006770521, 1.0079999e-06, -1.278912e-06, 0.011768455, 0.00069252035, 2.590826e-06, -1.271139e-06, 0.011418591, 0.00070671865, 4.188613e-06, -1.2580974e-06, 0.011061951, 0.0007196309, 5.7969696e-06, -1.2398594e-06, 0.010699177, 0.00073124404, 7.4115273e-06, -1.2165135e-06, 0.010330924, 0.00074154814, 9.02795e-06, -1.1881637e-06, 0.009957848, 0.0007505362, 1.0641949e-05, -1.154929e-06, 0.0095806075, 0.00075820443, 1.2249292e-05, -1.1169429e-06, 0.009199864, 0.0007645519, 1.3845814e-05, -1.0743521e-06, 0.008816276, 0.0007695808, 1.5427428e-05, -1.0273158e-06, 0.008430502, 0.00077329593, 1.699014e-05, -9.760051e-07, 0.008043197, 0.0007757053, 1.8530049e-05, -9.2060213e-07, 0.0076550124, 0.0007768197, 2.0043366e-05, -8.612991e-07, 0.0072665913, 0.0007766524, 2.1526417e-05, -7.982977e-07, 0.006878571, 0.0007752197, 2.2975652e-05, -7.318081e-07, 0.0064915796, 0.0007725403, 2.4387655e-05, -6.6204797e-07, 0.006106235, 0.0007686354, 2.5759146e-05, -5.892422e-07, 0.0057231444, 0.00076352886, 2.7086993e-05, -5.1362133e-07, 0.005342902, 0.0007572467, 2.8368218e-05, -4.3542153e-07, 0.004966089, 0.0007498172, 2.96e-05, -3.5488307e-07, 0.004593271, 0.00074127084, 3.0779676e-05, -2.7225e-07, 0.004224999, 0.0007316402, 3.1904754e-05, -1.8776915e-07, 0.003861806, 0.0007209598, 3.2972916e-05, -1.016894e-07, 0.003504208, 0.00070926594, 3.3982007e-05, -1.4260949e-08, 0.0031527025, 0.00069659663, 3.4930064e-05, 7.4265515e-08, 0.0028077674, 0.0006829916, 3.5815297e-05, 1.6363948e-07, 0.00246986, 0.0006684919, 3.663609e-05, 2.5361132e-07, 0.0021394175, 0.0006531401, 3.7391026e-05, 3.4393307e-07, 0.0018168548, 0.00063697994, 3.8078855e-05, 4.3435898e-07, 0.0015025649, 0.0006200564, 3.869852e-05, 5.246463e-07, 0.0011969181, 0.00060241536, 3.9249146e-05, 6.145557e-07, 0.0009002614, 0.0005841035, 3.973004e-05, 7.0385215e-07, 0.00061291846, 0.0005651685, 4.0140687e-05, 7.9230534e-07, 0.0003351888, 0.0005456585, 4.048076e-05, 8.796902e-07, 6.734773e-05, 0.0005256222, 4.0750107e-05, 9.657875e-07, -0.00019035382, 0.00050510874, 4.0948744e-05, 1.0503844e-06, -0.00043768962, 0.0004841674, 4.1076873e-05, 1.1332747e-06, -0.0006744581, 0.00046284776, 4.113486e-05, 1.2142597e-06, -0.0009004825, 0.00044119937, 4.112323e-05, 1.293148e-06, -0.0011156108, 0.00041927173, 4.1042673e-05, 1.3697564e-06, -0.0013197159, 0.00039711408, 4.0894043e-05, 1.4439103e-06, -0.0015126948, 0.0003747754, 4.0678347e-05, 1.5154434e-06, -0.0016944691, 0.00035230428, 4.0396728e-05, 1.5841987e-06, -0.0018649849, 0.00032974873, 4.005048e-05, 1.6500285e-06, -0.0020242117, 0.0003071562, 3.9641036e-05, 1.7127944e-06, -0.0021721425, 0.00028457335, 3.9169958e-05, 1.7723679e-06, -0.0023087943, 0.00026204612, 3.8638926e-05, 1.8286304e-06, -0.0024342055, 0.00023961939, 3.804975e-05, 1.8814732e-06, -0.0025484376, 0.00021733719, 3.7404352e-05, 1.9307977e-06, -0.0026515739, 0.00019524238, 3.670475e-05, 1.976516e-06, -0.0027437182, 0.00017337665, 3.5953068e-05, 2.0185496e-06, -0.0028249954, 0.00015178052, 3.5151523e-05, 2.0568316e-06, -0.00289555, 0.00013049312, 3.430242e-05, 2.0913042e-06, -0.0029555461, 0.000109552224, 3.3408134e-05, 2.1219207e-06, -0.003005166, 8.899417e-05, 3.2471118e-05, 2.1486442e-06, -0.00304461, 6.8853784e-05, 3.149389e-05, 2.1714486e-06, -0.003074095, 4.9164333e-05, 3.0479021e-05, 2.1903172e-06, -0.0030938545, 2.9957473e-05, 2.9429133e-05, 2.2052434e-06, -0.0031041377, 1.1263215e-05, 2.834689e-05, 2.216231e-06, -0.003105208, -6.8901313e-06, 2.7234997e-05, 2.2232928e-06, -0.0030973423, -2.447598e-05, 2.6096179e-05, 2.226451e-06, -0.0030808307, -4.1469506e-05, 2.4933186e-05, 2.2257375e-06, -0.0030559753, -5.7847665e-05, 2.3748784e-05, 2.2211932e-06, -0.0030230891, -7.3589224e-05, 2.2545744e-05, 2.2128672e-06, -0.0029824954, -8.8674766e-05, 2.1326836e-05, 2.2008176e-06, -0.0029345267, -0.00010308671, 2.0094829e-05, 2.1851106e-06, -0.0028795234, -0.00011680934, 1.8852472e-05, 2.16582e-06, -0.0028178345, -0.00012982874, 1.7602502e-05, 2.1430276e-06, -0.002749814, -0.00014213285, 1.6347625e-05, 2.1168223e-06, -0.0026758225, -0.00015371149, 1.5090519e-05, 2.0872997e-06, -0.002596225, -0.00016455624, 1.3833823e-05, 2.0545624e-06, -0.0025113896, -0.00017466056, 1.2580132e-05, 2.0187185e-06, -0.0024216885, -0.00018401962, 1.1331994e-05, 1.9798829e-06, -0.0023274948, -0.00019263044, 1.0091903e-05, 1.938175e-06, -0.002229183, -0.00020049176, 8.8622955e-06, 1.8937199e-06, -0.002127128, -0.00020760401, 7.64554e-06, 1.846647e-06, -0.0020217034, -0.00021396932, 6.443941e-06, 1.7970901e-06, -0.0019132824, -0.0002195915, 5.2597284e-06, 1.745187e-06, -0.0018022349, -0.0002244759, 4.0950563e-06, 1.6910788e-06, -0.0016889283, -0.00022862946, 2.9519979e-06, 1.6349095e-06, -0.001573726, -0.00023206066, 1.8325427e-06, 1.5768263e-06, -0.0014569864, -0.00023477942, 7.38593e-07, 1.5169782e-06, -0.0013390634, -0.0002367971, -3.2803908e-07, 1.4555162e-06, -0.001220304, -0.00023812639, -1.3656344e-06, 1.3925928e-06, -0.0011010494, -0.00023878133, -2.372569e-06, 1.3283615e-06, -0.0009816326, -0.00023877717, -3.3473168e-06, 1.2629763e-06, -0.0008623794, -0.00023813036, -4.288451e-06, 1.1965919e-06, -0.0007436065, -0.0002368585, -5.1946454e-06, 1.1293628e-06, -0.000625622, -0.00023498024, -6.0646767e-06, 1.0614427e-06, -0.0005087241, -0.00023251523, -6.897425e-06, 9.929848e-07, -0.00039320113, -0.00022948405, -7.691875e-06, 9.24141e-07, -0.00027933085, -0.00022590818, -8.447116e-06, 8.550617e-07, -0.00016738006, -0.00022180987, -9.162341e-06, 7.858955e-07, -5.7604266e-05, -0.0002172121, -9.83685e-06, 7.1678863e-07, 4.9752703e-05, -0.00021213855, -1.0470048e-05, 6.4788503e-07, 0.00015445899, -0.00020661348, -1.1061443e-05, 5.7932573e-07, 0.00025629502, -0.00020066166, -1.1610647e-05, 5.1124863e-07, 0.0003550537, -0.00019430835, -1.2117375e-05, 4.437883e-07, 0.00045054068, -0.0001875792, -1.2581445e-05, 3.7707576e-07, 0.00054257456, -0.00018050017, -1.3002771e-05, 3.11238e-07, 0.0006309869, -0.00017309746, -1.338137e-05, 2.46398e-07, 0.00071562245, -0.00016539752, -1.3717353e-05, 1.826743e-07, 0.00079633924, -0.00015742687, -1.4010926e-05, 1.2018099e-07, 0.00087300857, -0.0001492121, -1.4262389e-05, 5.9027336e-08, 0.00094551506, -0.0001407798, -1.447213e-05, -6.822579e-10, 0.0010137565, -0.0001321565, -1.4640624e-05, -5.8848492e-08, 0.0010776441, -0.00012336859, -1.4768433e-05, -1.153773e-07, 0.001137102, -0.00011444229, -1.4856199e-05, -1.7017996e-07, 0.0011920676, -0.000105403546, -1.4904645e-05, -2.2317325e-07, 0.0012424911, -9.627802e-05, -1.4914564e-05, -2.7427947e-07, 0.0012883353, -8.7091015e-05, -1.4886829e-05, -3.2342666e-07, 0.0013295759, -7.7867415e-05, -1.4822377e-05, -3.7054852e-07, 0.0013662007, -6.863166e-05, -1.4722211e-05, -4.1558457e-07, 0.0013982096, -5.940767e-05, -1.4587396e-05, -4.5848014e-07, 0.0014256142, -5.0218805e-05, -1.4419057e-05, -4.991864e-07, 0.001448438, -4.108784e-05, -1.4218371e-05, -5.3766047e-07, 0.0014667154, -3.203689e-05, -1.3986567e-05, -5.7386524e-07, 0.0014804917, -2.3087405e-05, -1.3724919e-05, -6.077694e-07, 0.0014898231, -1.4260112e-05, -1.34347465e-05, -6.3934755e-07, 0.0014947755, -5.5749824e-06, -1.3117407e-05, -6.6857996e-07, 0.001495425, 2.948796e-06, -1.27742915e-05, -6.9545274e-07, 0.0014918568, 1.1292848e-05, -1.2406825e-05, -7.199574e-07, 0.001484165, 1.9439643e-05, -1.2016456e-05, -7.4209134e-07, 0.0014724527, 2.7372516e-05, -1.1604659e-05, -7.6185705e-07, 0.0014568308, 3.507569e-05, -1.1172928e-05, -7.7926256e-07, 0.0014374178, 4.253429e-05, -1.072277e-05, -7.943212e-07, 0.0014143395, 4.973438e-05, -1.0255704e-05, -8.070512e-07, 0.0013877286, 5.666295e-05, -9.77326e-06, -8.1747595e-07, 0.0013577238, 6.330795e-05, -9.276969e-06, -8.2562354e-07, 0.0013244698, 6.965827e-05, -8.768362e-06, -8.3152685e-07, 0.0012881164, 7.570381e-05, -8.248969e-06, -8.3522303e-07, 0.0012488184, 8.143539e-05, -7.72031e-06, -8.3675377e-07, 0.0012067347, 8.684485e-05, -7.1838986e-06, -8.361648e-07, 0.0011620284, 9.1924965e-05, -6.641231e-06, -8.33506e-07, 0.0011148656, 9.66695e-05, -6.093788e-06, -8.288307e-07, 0.0010654157, 0.000101073194, -5.543032e-06, -8.221961e-07, 0.00101385, 0.000105131716, -4.9903992e-06, -8.1366267e-07, 0.00096034206, 0.00010884172, -4.4373014e-06, -8.032939e-07, 0.0009050668, 0.00011220076, -3.8851213e-06, -7.9115654e-07, 0.00084820006, 0.000115207346, -3.3352094e-06, -7.7731977e-07, 0.0007899183, 0.00011786087, -2.7888827e-06, -7.618556e-07, 0.000730398, 0.00012016164, -2.2474212e-06, -7.448381e-07, 0.0006698153, 0.00012211081, -1.7120661e-06, -7.263435e-07, 0.0006083455, 0.00012371042, -1.1840173e-06, -7.0645007e-07, 0.0005461627, 0.0001249633, -6.6443147e-07, -6.8523747e-07, 0.0004834394, 0.0001258731, -1.544205e-07, -6.6278704e-07, 0.00042034604, 0.00012644428, 3.4495065e-07, -6.391811e-07, 0.0003570507, 0.000126682, 8.3266536e-07, -6.145032e-07, 0.00029371865, 0.00012659217, 1.3077569e-06, -5.888375e-07, 0.00023051204, 0.0001261814, 1.7693094e-06, -5.622688e-07, 0.00016758955, 0.00012545697, 2.2164597e-06, -5.348822e-07, 0.00010510606, 0.00012442676, 2.6483974e-06, -5.0676306e-07, 4.3212363e-05, 0.00012309928, 3.0643669e-06, -4.7799654e-07, -1.7945164e-05, 0.000121483616, 3.4636669e-06, -4.4866758e-07, -7.8224795e-05, 0.00011958936, 3.8456515e-06, -4.188608e-07, -0.00013748975, 0.00011742662, 4.2097313e-06, -3.8866e-07, -0.0001956084, 0.00011500597, 4.555372e-06, -3.5814827e-07, -0.00025245454, 0.0001123384, 4.8820966e-06, -3.274076e-07, -0.00030790752, 0.000109435314, 5.189484e-06, -2.9651886e-07, -0.00036185252, 0.000106308464, 5.4771685e-06, -2.6556154e-07, -0.0004141807, 0.00010296991, 5.7448415e-06, -2.3461364e-07, -0.0004647892, 9.943203e-05, 5.9922486e-06, -2.0375144e-07, -0.00051358156, 9.5707415e-05, 6.219192e-06, -1.7304944e-07, -0.0005604676, 9.1808906e-05, 6.425527e-06, -1.425802e-07, -0.00060536363, 8.774949e-05, 6.611162e-06, -1.1241415e-07, -0.0006481924, 8.354231e-05, 6.7760593e-06, -8.2619515e-08, -0.0006888835, 7.9200625e-05, 6.9202333e-06, -5.326218e-08, -0.0007273728, 7.473775e-05, 7.043747e-06, -2.4405603e-08, -0.00076360325, 7.016705e-05, 7.1467143e-06, 3.889324e-09, -0.0007975241, 6.5501896e-05, 7.2292974e-06, 3.1564344e-08, -0.0008290916, 6.075562e-05, 7.291704e-06, 5.856393e-08, -0.0008582684, 5.5941502e-05, 7.3341894e-06, 8.483536e-08, -0.00088502397, 5.107273e-05, 7.3570504e-06, 1.1032878e-07, -0.0009093342, 4.616237e-05, 7.3606266e-06, 1.3499728e-07, -0.00093118154, 4.1223335e-05, 7.3452993e-06, 1.5879695e-07, -0.00095055485, 3.6268357e-05, 7.311487e-06, 1.8168689e-07, -0.00096744933, 3.130996e-05, 7.2596463e-06, 2.0362927e-07, -0.0009818663, 2.6360438e-05, 7.1902678e-06, 2.245894e-07, -0.0009938133, 2.1431819e-05, 7.1038767e-06, 2.4453567e-07, -0.0010033036, 1.653585e-05, 7.001028e-06, 2.634396e-07, -0.0010103564, 1.1683969e-05, 6.882307e-06, 2.8127587e-07, -0.0010149967, 6.887285e-06, 6.7483256e-06, 2.9802231e-07, -0.0010172547, 2.1565565e-06, 6.5997215e-06, 3.1365983e-07, -0.001017166, -2.4978276e-06, 6.437155e-06, 3.2817246e-07, -0.0010147712, -7.0658666e-06, 6.261308e-06, 3.4154735e-07, -0.0010101161, -1.1537964e-05, 6.0728808e-06, 3.5377462e-07, -0.0010032507, -1.5904945e-05, 5.872591e-06, 3.6484752e-07, -0.00099423, -2.0158068e-05, 5.6611707e-06, 3.7476218e-07, -0.0009831131, -2.4289038e-05, 5.4393654e-06, 3.8351766e-07, -0.0009699627, -2.8290024e-05, 5.2079304e-06, 3.9111592e-07, -0.0009548459, -3.2153654e-05, 4.9676296e-06, 3.9756165e-07, -0.0009378331, -3.5873047e-05, 4.7192348e-06, 4.0286236e-07, -0.000918998, -3.94418e-05, 4.463521e-06, 4.0702812e-07, -0.0008984174, -4.2853997e-05, 4.2012653e-06, 4.1007166e-07, -0.00087617093, -4.610423e-05, 3.933247e-06, 4.1200818e-07, -0.00085234095, -4.918758e-05, 3.660244e-06, 4.1285523e-07, -0.00082701194, -5.2099636e-05, 3.383029e-06, 4.1263277e-07, -0.0008002705, -5.4836495e-05, 3.1023721e-06, 4.113629e-07, -0.0007722052, -5.7394747e-05, 2.8190354e-06, 4.090699e-07, -0.000742906, -5.9771486e-05, 2.5337724e-06, 4.0578007e-07, -0.0007124644, -6.196431e-05, 2.2473273e-06, 4.015216e-07, -0.0006809727, -6.397131e-05, 1.9604315e-06, 3.9632445e-07, -0.00064852426, -6.5791064e-05, 1.6738037e-06, 3.9022038e-07, -0.000615213, -6.742264e-05, 1.3881476e-06, 3.8324262e-07, -0.00058113306, -6.8865564e-05, 1.1041507e-06, 3.7542603e-07, -0.0005463789, -7.011986e-05, 8.224829e-07, 3.6680666e-07, -0.0005110446, -7.118599e-05, 5.437951e-07, 3.574219e-07, -0.0004752241, -7.206488e-05, 2.6871828e-07, 3.4731028e-07, -0.0004390107, -7.275787e-05, -2.1380147e-09, 3.365113e-07, -0.00040249692, -7.326677e-05, -2.6818645e-07, 3.250654e-07, -0.00036577426, -7.359374e-05, -5.2886304e-07, 3.1301374e-07, -0.00032893306, -7.3741416e-05, -7.8362797e-07, 3.003982e-07, -0.00029206224, -7.3712756e-05, -1.0319665e-06, 2.8726117e-07, -0.00025524915, -7.351113e-05, -1.2733898e-06, 2.7364553e-07, -0.00021857933, -7.314025e-05, -1.5074353e-06, 2.5959437e-07, -0.00018213644, -7.2604154e-05, -1.7336679e-06, 2.4515114e-07, -0.000146002, -7.1907234e-05, -1.95168e-06, 2.303593e-07, -0.00011025524, -7.105417e-05, -2.1610917e-06, 2.1526229e-07, -7.497303e-05, -7.004994e-05, -2.361552e-06, 1.9990347e-07, -4.022964e-05, -6.889978e-05, -2.552739e-06, 1.8432597e-07, -6.096666e-06, -6.7609195e-05, -2.7343588e-06, 1.6857263e-07, 2.7357097e-05, -6.618392e-05, -2.9061473e-06, 1.5268581e-07, 6.0065784e-05, -6.462991e-05, -3.0678696e-06, 1.3670744e-07, 9.196656e-05, -6.295331e-05, -3.2193198e-06, 1.2067878e-07, 0.0001229997, -6.116045e-05, -3.360321e-06, 1.0464043e-07, 0.0001531087, -5.925783e-05, -3.4907257e-06, 8.86322e-08, 0.00018224033, -5.7252073e-05, -3.6104145e-06, 7.2693055e-08, 0.0002103447, -5.514994e-05, -3.7192976e-06, 5.686101e-08, 0.00023737534, -5.295829e-05, -3.817312e-06, 4.1173067e-08, 0.00026328923, -5.0684073e-05, -3.904424e-06, 2.5665162e-08, 0.0002880468, -4.8334296e-05, -3.9806255e-06, 1.037207e-08, 0.0003116121, -4.591602e-05, -4.0459363e-06, -4.67264e-09, 0.00033395257, -4.343634e-05, -4.1004023e-06, -1.9436667e-08, 0.00035503937, -4.090236e-05, -4.1440944e-06, -3.388903e-08, 0.00037484706, -3.832118e-05, -4.1771095e-06, -4.800012e-08, 0.00039335384, -3.5699883e-05, -4.1995677e-06, -6.1741744e-08, 0.00041054143, -3.30455e-05, -4.211613e-06, -7.508717e-08, 0.00042639498, -3.0365021e-05, -4.213412e-06, -8.801115e-08, 0.00044090324, -2.7665357e-05, -4.2051524e-06, -1.0048996e-07, 0.0004540583, -2.4953339e-05, -4.187044e-06, -1.1250146e-07, 0.0004658556, -2.2235692e-05, -4.1593153e-06, -1.2402504e-07, 0.00047629414, -1.9519026e-05, -4.1222147e-06, -1.350417e-07, 0.0004853759, -1.6809823e-05, -4.0760087e-06, -1.4553409e-07, 0.00049310626, -1.4114422e-05, -4.02098e-06, -1.5548643e-07, 0.0004994936, -1.1439008e-05, -3.9574284e-06, -1.648846e-07, 0.0005045496, -8.789597e-06, -3.8856674e-06, -1.7371607e-07, 0.0005082885, -6.172028e-06, -3.8060255e-06, -1.8197001e-07, 0.00051072787, -3.5919504e-06, -3.7188438e-06, -1.8963712e-07, 0.00051188766, -1.054814e-06, -3.624475e-06, -1.9670982e-07, 0.0005117907, 1.4341393e-06, -3.5232827e-06, -2.0318203e-07, 0.0005104623, 3.8698854e-06, -3.4156399e-06, -2.0904932e-07, 0.00050793047, 6.2476247e-06, -3.3019278e-06, -2.143088e-07, 0.00050422514, 8.562791e-06, -3.182536e-06, -2.1895912e-07, 0.00049937883, 1.0811055e-05, -3.0578592e-06, -2.2300044e-07, 0.00049342593, 1.2988336e-05, -2.928298e-06, -2.2643444e-07, 0.00048640295, 1.5090798e-05, -2.7942576e-06, -2.2926419e-07, 0.0004783482, 1.7114864e-05, -2.6561452e-06, -2.3149421e-07, 0.0004693017, 1.9057215e-05, -2.5143706e-06, -2.331304e-07, 0.0004593051, 2.091479e-05, -2.369345e-06, -2.3417998e-07, 0.0004484015, 2.2684793e-05, -2.221479e-06, -2.3465147e-07, 0.00043663534, 2.4364694e-05, -2.0711823e-06, -2.3455462e-07, 0.0004240522, 2.5952228e-05, -1.9188628e-06, -2.3390038e-07, 0.00041069882, 2.7445398e-05, -1.7649253e-06, -2.3270088e-07, 0.0003966228, 2.8842473e-05, -1.6097708e-06, -2.309693e-07, 0.0003818726, 3.0141984e-05, -1.4537956e-06, -2.2871988e-07, 0.0003664973, 3.134273e-05, -1.2973902e-06, -2.2596784e-07, 0.0003505465, 3.244377e-05, -1.1409387e-06, -2.2272935e-07, 0.00033407027, 3.344442e-05, -9.84818e-07, -2.1902143e-07, 0.0003171189, 3.434425e-05, -8.293968e-07, -2.1486191e-07, 0.00029974285, 3.514309e-05, -6.750352e-07, -2.102694e-07, 0.00028199263, 3.5841003e-05, -5.2208367e-07, -2.0526318e-07, 0.00026391863, 3.6438305e-05, -3.7088242e-07, -1.998632e-07, 0.000245571, 3.6935544e-05, -2.2176111e-07, -1.940899e-07, 0.00022699962, 3.7333502e-05, -7.5037846e-08, -1.8796436e-07, 0.00020825388, 3.7633177e-05, 6.8981144e-08, -1.81508e-07, 0.00018938263, 3.7835795e-05, 2.1000207e-07, -1.7474268e-07};
endpackage
`endif
