`ifndef COEFFICIENTS_SV_
`define COEFFICIENTS_SV_
package Coefficients;
	localparam real Lfr[0:2] = {0.9616946545986035, 0.9293198051200361, 0.9616946545986016};
	localparam real Lfi[0:2] = {0.061059134464848674, 2.110941629829277e-15, -0.06105913446485091};
	localparam real Lbr[0:2] = {0.9616946545986075, 0.9293198051200214, 0.9616946545986091};
	localparam real Lbi[0:2] = {0.06105913446485922, -3.198835171898916e-15, -0.0610591344648556};
	localparam real Wfr[0:2] = {1.1135647654883724e-05, -0.0005307564331930271, 1.1135647654962437e-05};
	localparam real Wfi[0:2] = {-0.0009207389130005212, -7.544389062598468e-18, 0.0009207389130004935};
	localparam real Wbr[0:2] = {-1.1269258956132365e-05, 0.000533843812413026, -1.1269258956024108e-05};
	localparam real Wbi[0:2] = {0.0009233839399884489, -1.4503522108469972e-17, -0.000923383939988464};
	localparam real Ffr[0:2][0:59] = '{
		'{11.182709042544154, -1.5872948617600278, -0.0270186711577089, 10.335170870306293, -1.586267003551229, -0.01006330868911368, 9.49446322365076, -1.577071072215828, 0.00573346772374899, 8.66446621060493, -1.5603381697337786, 0.02037232627843925, 7.84872719332538, -1.5366934862923367, 0.033859903435438515, 7.050466120820197, -1.506753474291275, 0.04620834321377214, 6.272582181914673, -1.471123269564328, 0.05743484077329894, 5.5176616496094635, -1.4303943555599736, 0.06756119234886054, 4.7879867909920915, -1.3851424652663495, 0.07661335342099651, 4.08554572031364, -1.3359257148023622, 0.0846210068305411, 3.412043076682403, -1.2832829618274568, 0.09161714237082573, 2.768911412008245, -1.227732381243499, 0.0976376492220481, 2.1573231793086967, -1.169770250070782, 0.10272092242819648, 1.5782032162164334, -1.1098699328731503, 0.10690748445823406, 1.032241623464902, -1.048481058681225, 0.11023962274048313, 0.5199069432343384, -0.9860288800141805, 0.11276104391267754, 0.0414595474752244, -0.9229138043256777, 0.11451654539027972, -0.4030348483456594, -0.8595110879946404, 0.11555170472264954, -0.8136916252445383, -0.7961706828425748, 0.11591258708069618, -1.1907937282198289, -0.733217225082154, 0.1156454711009044},
		'{-21.938581601088295, 2.995512590835637, -0.4181464982722033, -20.387958378133384, 2.7837891771499885, -0.38859182228594946, -18.946933506762324, 2.587030415604293, -0.36112607655801826, -17.607760554126646, 2.404178601668988, -0.3356016150906608, -16.36324060676123, 2.2342507895767842, -0.31188122753402225, -15.20668357180761, 2.0763335083587844, -0.2898374015925152, -14.131872213474303, 1.9295778513521862, -0.26935163756445385, -13.133028731407192, 1.7931949127825517, -0.25031381133016084, -12.204783701307166, 1.6664515468893208, -0.23262158236419855, -11.34214721083097, 1.5486664267971664, -0.21617984358941142, -10.540482035612197, 1.4392063819470853, -0.20090021011539172, -9.795478711206368, 1.3374829943985778, -0.18670054411301015, -9.103132366955764, 1.2429494357058484, -0.17350451327090727, -8.459721197241224, 1.155097527364218, -0.16124118046036628, -7.861786454390052, 1.0734550090247506, -0.14984462240275215, -7.306113855689103, 0.9975829997920078, -0.13925357528961102, -6.789716304553792, 0.9270736389577696, -0.1294111054504096, -6.309817832968262, 0.8615478934881572, -0.12026430329754308, -5.863838678876994, 0.8006535204779919, -0.11176399890336965, -5.449381418309298, 0.7440631736192782, -0.10386449768031542},
		'{11.182709042544008, -1.5872948617599003, -0.02701867115773409, 10.335170870306213, -1.5862670035511124, -0.010063308689137435, 9.494463223650737, -1.5770710722157222, 0.005733467723726644, 8.66446621060496, -1.560338169733682, 0.02037232627841827, 7.848727193325459, -1.5366934862922486, 0.03385990343541885, 7.050466120820317, -1.506753474291195, 0.04620834321375375, 6.272582181914835, -1.4711232695642555, 0.05743484077328178, 5.51766164960966, -1.4303943555599075, 0.06756119234884456, 4.787986790992321, -1.3851424652662896, 0.0766133534209816, 4.085545720313899, -1.335925714802308, 0.08462100683052722, 3.412043076682689, -1.2832829618274075, 0.09161714237081282, 2.7689114120085536, -1.227732381243454, 0.09763764922203609, 2.1573231793090297, -1.1697702500707416, 0.10272092242818534, 1.5782032162167852, -1.1098699328731136, 0.1069074844582237, 1.0322416234652705, -1.0484810586811917, 0.11023962274047351, 0.5199069432347234, -0.9860288800141503, 0.11276104391266856, 0.04145954747562364, -0.9229138043256506, 0.11451654539027137, -0.4030348483452477, -0.8595110879946157, 0.11555170472264173, -0.8136916252441151, -0.7961706828425524, 0.11591258708068888, -1.190793728219396, -0.733217225082134, 0.11564547110089755}};
localparam real Ffi[0:2][0:59] = '{
	'{6.865158563313831, 0.9789529486238033, -0.2607374486577057, 7.284992828420722, 0.8445349673954841, -0.25239954730307346, 7.63699524976859, 0.7153286734988558, -0.243345752382883, 7.924181215541831, 0.59163316692591, -0.2336742287091997, 8.149687524476708, 0.4736975559994802, -0.22347934005749184, 8.316747418013342, 0.36172323329034184, -0.21285143034968224, 8.428666894461188, 0.25586623690731647, -0.20187664134926878, 8.48880233668288, 0.15623967879533007, -0.19063676520816716, 8.500539475727102, 0.0629162226397747, -0.17920913014242879, 8.467273704298275, -0.024069405039462977, -0.16766651746490363, 8.392391745945885, -0.10471788602098675, -0.15607710816654435, 8.279254678392606, -0.17906277814992066, -0.1445044572136683, 8.131182302497713, -0.2471679931375501, -0.1330074937153766, 7.951438841968359, -0.3091252967802977, -0.12164054511273849, 7.743219953080495, -0.3650518429846133, -0.11045338354854686, 7.509641018346121, -0.4150877519955354, -0.0994912925927015, 7.25372669325403, -0.459393742254467, -0.08879515252284575, 6.978401670905746, -0.4981488243599561, -0.07840154239205344, 6.686482625552862, -0.5315480646774414, -0.06834285715442086, 6.380671292701894, -0.5598004252431834, -0.05864743816467374},
	'{-1.511614781428562e-12, 1.1297547625164232e-13, 2.4565125697653787e-15, -1.4510846192949011e-12, 1.1131369980419221e-13, 1.400202932039151e-15, -1.3915594657034476e-12, 1.093224422719362e-13, 4.809416612564959e-16, -1.3331996421775012e-12, 1.0705658094933578e-13, -3.153674577102424e-16, -1.276137786416269e-12, 1.045648816404619e-13, -1.001512644673301e-15, -1.2204819647744066e-12, 1.0189058843171027e-13, -1.5890886025368682e-15, -1.1663184830600398e-12, 9.907196062512682e-14, -2.0886013473312195e-15, -1.113714422748103e-12, 9.61427613554186e-14, -2.509564181872787e-15, -1.0627199273825119e-12, 9.313270203831053e-14, -2.860585541292309e-15, -1.0133702618104461e-12, 9.006784645296719e-14, -3.1494493799723083e-15, -9.65687664939119e-13, 8.69709779442979e-14, -3.383188715394155e-15, -9.19683014915486e-13, 8.386193293986196e-14, -3.56815289464843e-15, -8.753573239890588e-13, 8.075790370872673e-14, -3.710069103573102e-15, -8.327030788151616e-13, 7.767371304410085e-14, -3.814098596341246e-15, -7.917054405793657e-13, 7.462206332611939e-14, -3.8848880845370525e-15, -7.523433180630883e-13, 7.161376221418339e-14, -3.926616689071143e-15, -7.145903256159972e-13, 6.865792702826842e-14, -3.943038825450081e-15, -6.784156369441348e-13, 6.576216970424933e-14, -3.937523362705501e-15, -6.437847446555604e-13, 6.29327640482796e-14, -3.9130893684982636e-15, -6.106601346204022e-13, 6.017479686845878e-14, -3.872438727351409e-15},
	'{-6.865158563312287, -0.9789529486239181, 0.2607374486577031, -7.28499282841924, -0.8445349673955967, 0.25239954730307207, -7.636995249767168, -0.7153286734989662, 0.24334575238288267, -7.92418121554047, -0.5916331669260178, 0.23367422870920027, -8.149687524475404, -0.4736975559995853, 0.2234793400574932, -8.316747418012099, -0.36172323329044404, 0.2128514303496843, -8.42866689446, -0.2558662369074155, 0.20187664134927133, -8.488802336681744, -0.156239678795426, 0.1906367652081702, -8.500539475726018, -0.06291622263986762, 0.17920913014243214, -8.467273704297241, 0.02406940503937338, 0.16766651746490727, -8.392391745944899, 0.10471788602090015, 0.15607710816654818, -8.279254678391666, 0.17906277814983712, 0.14450445721367225, -8.131182302496823, 0.24716799313746934, 0.13300749371538073, -7.951438841967512, 0.30912529678021977, 0.12164054511274267, -7.743219953079692, 0.36505184298453813, 0.11045338354855103, -7.5096410183453575, 0.4150877519954625, 0.09949129259270564, -7.2537266932533075, 0.45939374225439655, 0.08879515252284988, -6.978401670905061, 0.49814882435988783, 0.07840154239205747, -6.686482625552214, 0.5315480646773754, 0.06834285715442481, -6.380671292701284, 0.5598004252431192, 0.05864743816467761}};
	localparam real Fbr[0:2][0:59] = '{
		'{-11.151414532990982, -1.805772860263286, -0.03939046885537871, -10.306351328017413, -1.7878609332011912, -0.05602552426643666, -9.468091630842856, -1.7619393269508046, -0.0711815027250545, -8.640504760610268, -1.7287147302963524, -0.084885289618672, -7.827128257507071, -1.6888813065336126, -0.09716939519664919, -7.031173197465227, -1.6431179814423722, -0.10807138396221096, -6.255530823461821, -1.5920860041055795, -0.1176333185550012, -5.502780364941836, -1.5364267737626065, -0.12590121997871473, -4.77519791988723, -1.4767599249883687, -0.13292454581091726, -4.0747662774962885, -1.413681662698405, -0.13875568782182224, -3.403185563265524, -1.3477633377890572, -0.14344949022606096, -2.7618845924353717, -1.2795502536280468, -0.14706278959686842, -2.1520328222247596, -1.2095606931101193, -0.1496539772860436, -1.5745527979938627, -1.138285155581014, -0.1512825850158852, -1.0301329933968657, -1.066185792606558, -0.15200889414133617, -0.5192409496765902, -0.9936960313177863, -0.1518935689220108, -0.042136624472310036, -0.9212203738932379, -0.15099731399477548, 0.40111413417563657, -0.8491343616413537, -0.14938055609820386, 0.8106260675698196, -0.7777846921146381, -0.14710314997056073, 1.1866810133960417, -0.7074894777183283, -0.1442241082229698},
		'{21.811704189790145, 3.414218810004178, 0.5463712179502375, 20.270048686991334, 3.1729011591501943, 0.5077535937887034, 18.83735769556813, 2.948639886886548, 0.4718654708287084, 17.505929582621512, 2.740229445050529, 0.43851392739340245, 16.26860706816664, 2.5465494938585023, 0.407519677547652, 15.118738750162827, 2.366558879361073, 0.3787161073211579, 14.050143348961832, 2.1992900365728882, 0.35194837905151155, 13.057076478965577, 2.0438437881903213, 0.32707259903245817, 12.134199768869506, 1.8993845109367957, 0.30395504399294293, 11.276552164493216, 1.76513564355177, 0.28247144224876924, 10.479523259932591, 1.6403755122759345, 0.26250630566259764, 9.738828513671288, 1.5244334513919269, 0.243952308821142, 9.05048621642231, 1.4166861979659873, 0.226709712092243, 8.410796086887022, 1.3165545414099753, 0.21068582546037942, 7.816319380370085, 1.2235002098529972, 0.19579451025839065, 7.263860403321375, 1.137022976584893, 0.18195571611689765, 6.75044933443366, 1.0566579710168593, 0.16909505064222927, 6.273326259948468, 0.9819731797039051, 0.15714337950959667, 5.829926337349622, 0.9125671239955208, 0.14603645482175992, 5.417866007689831, 0.8480667018304557, 0.13571456973537674},
		'{-11.151414532991534, -1.805772860263508, -0.03939046885542044, -10.306351328017865, -1.787860933201394, -0.056025524266475876, -9.46809163084321, -1.7619393269509898, -0.07118150272509124, -8.640504760610536, -1.7287147302965211, -0.08488528961870637, -7.827128257507262, -1.6888813065337662, -0.09716939519668126, -7.031173197465346, -1.6431179814425116, -0.10807138396224081, -6.255530823461873, -1.5920860041057059, -0.11763331855502893, -5.502780364941829, -1.5364267737627206, -0.12590121997874043, -4.775197919887169, -1.4767599249884724, -0.13292454581094104, -4.0747662774961775, -1.4136816626984983, -0.13875568782184422, -3.403185563265366, -1.3477633377891414, -0.14344949022608125, -2.7618845924351745, -1.279550253628123, -0.14706278959688712, -2.152032822224525, -1.2095606931101877, -0.1496539772860608, -1.5745527979935945, -1.1382851555810758, -0.15128258501590106, -1.030132993396565, -1.0661857926066132, -0.15200889414135074, -0.5192409496762616, -0.9936960313178353, -0.15189356892202424, -0.042136624471956985, -0.9212203738932818, -0.15099731399478786, 0.40111413417601405, -0.8491343616413929, -0.1493805560982153, 0.810626067570217, -0.7777846921146729, -0.14710314997057128, 1.186681013396458, -0.7074894777183593, -0.14422410822297957}};
localparam real Fbi[0:2][0:59] = '{
	'{-6.844257181761263, 0.839494803128127, 0.2971532610985211, -7.262981265841217, 0.6970787368438206, 0.2833655548605176, -7.614067151388824, 0.5612116539322515, 0.2690902693870797, -7.900521159258719, 0.43213175740187704, 0.254436392727754, -8.125470709424661, 0.3100249760071395, 0.239507096508718, -8.292139424100077, 0.19502773142730456, 0.22439961528368566, -8.403823509053161, 0.08722976504161395, 0.2092051653471524, -8.463869444545367, -0.013322994641890462, 0.19400890061357687, -8.475653008273333, -0.10662554170493277, 0.1788899031446592, -8.442559644175782, -0.19271089633349503, 0.16392120589953224, -8.36796618298429, -0.2716472176200362, 0.1491698452884612, -8.255223912954202, -0.34353493999064305, 0.13469694112858582, -8.107642992308591, -0.4085039464476744, 0.12055780162937184, -7.9284781885620434, -0.46671079068518334, 0.10680205107481665, -7.720915924056495, -0.5183359790194046, 0.09347377791814221, -7.488062601730906, -0.5635813219843838, 0.08061170106178434, -7.232934180350318, -0.6026673643774283, 0.06824935216006245, -6.9584469641260105, -0.635830901504119, 0.05641527185311042, -6.667409567853507, -0.6633225883713167, 0.04513321791762789, -6.362516015363863, -0.6854046476117446, 0.034422383401960015},
	'{-2.0079275152704267e-12, -1.6700790873444264e-13, 1.6408940462268885e-15, -1.9357788537075974e-12, -1.661252804125948e-13, -2.228361336302923e-16, -1.8637981717590542e-12, -1.6453310104338997e-13, -1.8313060867483817e-15, -1.7923221561044005e-12, -1.6233608237687268e-13, -3.21128888014363e-15, -1.7216390600889137e-12, -1.5962767876632377e-13, -4.387048130592713e-15, -1.6519938682963006e-12, -1.5649115541081735e-13, -5.380558991554908e-15, -1.5835929730133602e-12, -1.5300056182905765e-13, -6.211710437732151e-15, -1.5166084057850922e-12, -1.4922161862442982e-13, -6.898490387058031e-15, -1.4511816635906775e-12, -1.4521252493527962e-13, -7.45715507567253e-15, -1.3874271658053443e-12, -1.4102469335238494e-13, -7.902383987074482e-15, -1.3254353750259799e-12, -1.36703418523115e-13, -8.247421531374013e-15, -1.2652756120069312e-12, -1.322884851449319e-13, -8.504206573677931e-15, -1.206998592356021e-12, -1.2781472057604274e-13, -8.683490821473794e-15, -1.1506387102603157e-12, -1.2331249685479535e-13, -8.794946998825265e-15, -1.0962160923290733e-12, -1.1880818651874717e-13, -8.84726765969243e-15, -1.0437384426414088e-12, -1.1432457624636875e-13, -8.848255423229301e-15, -9.932026982536971e-13, -1.0988124200646139e-13, -8.804905350010414e-15, -9.445965127429133e-13, -1.0549488909014669e-13, -8.723480119360304e-15, -8.978995838244162e-13, -1.0117966011551167e-13, -8.609578613898657e-15, -8.530848396745484e-13, -9.69474138336128e-14, -8.468198467697074e-15},
	'{6.844257181763314, -0.8394948031279555, -0.2971532610985227, 7.262981265843196, -0.6970787368436502, -0.2833655548605173, 7.614067151390728, -0.5612116539320828, -0.2690902693870776, 7.90052115926055, -0.4321317574017109, -0.2544363927277505, 8.125470709426423, -0.3100249760069765, -0.23950709650871327, 8.292139424101766, -0.1950277314271452, -0.2243996152836799, 8.403823509054783, -0.08722976504145807, -0.2092051653471458, 8.46386944454692, 0.013322994642042008, -0.19400890061356962, 8.475653008274822, 0.10662554170507998, -0.17888990314465145, 8.442559644177207, 0.1927108963336377, -0.1639212058995241, 8.367966182985654, 0.2716472176201744, -0.1491698452884528, 8.255223912955504, 0.3435349399907765, -0.13469694112857733, 8.107642992309836, 0.40850394644780336, -0.1205578016293633, 7.928478188563233, 0.4667107906853079, -0.10680205107480815, 7.720915924057629, 0.518335979019525, -0.09347377791813374, 7.488062601731988, 0.5635813219844998, -0.08061170106177601, 7.23293418035135, 0.6026673643775402, -0.06824935216005434, 6.958446964126994, 0.635830901504227, -0.05641527185310252, 6.667409567854442, 0.6633225883714209, -0.04513321791762025, 6.362516015364752, 0.6854046476118452, -0.034422383401952625}};
	localparam real hf[0:1199] = {0.024535134, 0.00017748146, -0.00025881003, 0.024466371, 4.235018e-05, -0.0002587647, 0.024331018, -9.094456e-05, -0.00025631813, 0.024130605, -0.00022130465, -0.00025172948, 0.023867166, -0.0003477636, -0.00024524517, 0.023543173, -0.00046947942, -0.000237099, 0.023161484, -0.0005857277, -0.0002275121, 0.022725265, -0.0006958946, -0.00021669304, 0.022237957, -0.00079946994, -0.00020483795, 0.021703204, -0.00089604076, -0.00019213071, 0.021124823, -0.0009852841, -0.00017874302, 0.020506745, -0.001066961, -0.00016483472, 0.019852985, -0.0011409101, -0.00015055398, 0.019167598, -0.0012070411, -0.0001360376, 0.01845465, -0.0012653291, -0.00012141128, 0.017718183, -0.0013158086, -0.00010678994, 0.016962186, -0.0013585682, -9.22781e-05, 0.016190572, -0.0013937445, -7.7970166e-05, 0.015407158, -0.0014215177, -6.395087e-05, 0.014615638, -0.0014421061, -5.029563e-05, 0.013819575, -0.0014557614, -3.7070942e-05, 0.013022378, -0.0014627642, -2.4334788e-05, 0.012227292, -0.0014634201, -1.2137063e-05, 0.011437392, -0.001458055, -5.1998336e-07, 0.010655567, -0.0014470116, 1.0481489e-05, 0.009884519, -0.0014306457, 2.0839223e-05, 0.0091267545, -0.0014093232, 3.0531493e-05, 0.008384588, -0.0013834162, 3.9542574e-05, 0.00766013, -0.0013533011, 4.7862304e-05, 0.0069552967, -0.0013193549, 5.548569e-05, 0.006271805, -0.0012819533, 6.2412495e-05, 0.005611177, -0.0012414687, 6.864687e-05, 0.004974743, -0.0011982674, 7.419692e-05, 0.0043636453, -0.0011527084, 7.907438e-05, 0.0037788455, -0.0011051416, 8.329421e-05, 0.0032211267, -0.0010559057, 8.687428e-05, 0.0026911027, -0.0010053284, 8.983501e-05, 0.0021892241, -0.00095372356, 9.219905e-05, 0.0017157864, -0.0009013915, 9.399097e-05, 0.0012709373, -0.00084861775, 9.523697e-05, 0.0008546855, -0.00079567236, 9.596458e-05, 0.0004669088, -0.00074280956, 9.620242e-05, 0.00010736289, -0.0006902673, 9.5979936e-05, -0.00022430973, -0.00063826714, 9.5327174e-05, -0.0005285711, -0.0005870139, 9.427453e-05, -0.00080597884, -0.0005366958, 9.28526e-05, -0.0010571777, -0.00048748465, 9.109192e-05, -0.0012828903, -0.00043953562, 8.902286e-05, -0.0014839094, -0.00039298795, 8.6675434e-05, -0.0016610889, -0.0003479649, 8.407914e-05, -0.0018153363, -0.00030457444, 8.126284e-05, -0.0019476044, -0.0002629095, 7.825468e-05, -0.002058884, -0.00022304854, 7.50819e-05, -0.0021501961, -0.00018505605, 7.177084e-05, -0.0022225862, -0.00014898326, 6.8346795e-05, -0.0022771163, -0.0001148686, 6.4833956e-05, -0.0023148593, -8.273844e-05, 6.1255385e-05, -0.0023368932, -5.260775e-05, 5.7632937e-05, -0.002344295, -2.4480756e-05, 5.398723e-05, -0.0023381358, 1.6483531e-06, 5.0337643e-05, -0.0023194766, 2.579473e-05, 4.6702255e-05, -0.0022893632, 4.798216e-05, 4.3097876e-05, -0.0022488215, 6.824238e-05, 3.9540028e-05, -0.0021988559, 8.6614345e-05, 3.604295e-05, -0.0021404433, 0.000103143604, 3.2619617e-05, -0.0020745327, 0.00011788157, 2.9281751e-05, -0.0020020404, 0.0001308849, 2.603985e-05, -0.0019238496, 0.00014221483, 2.2903216e-05, -0.0018408066, 0.00015193659, 1.9879992e-05, -0.0017537207, 0.00016011875, 1.6977188e-05, -0.001663362, 0.00016683273, 1.4200738e-05, -0.0015704606, 0.00017215217, 1.1555529e-05, -0.0014757058, 0.0001761524, 9.045456e-06, -0.0013797453, 0.00017891006, 6.673466e-06, -0.0012831856, 0.00018050248, 4.44161e-06, -0.0011865911, 0.00018100737, 2.351094e-06, -0.0010904848, 0.00018050229, 4.0232976e-07, -0.0009953484, 0.00017906439, -1.4050113e-06, -0.0009016233, 0.00017676991, -3.071946e-06, -0.0008097103, 0.00017369405, -4.6001255e-06, -0.00071997166, 0.00016991043, -5.9917847e-06, -0.0006327311, 0.00016549104, -7.2496896e-06, -0.00054827565, 0.00016050591, -8.377085e-06, -0.0004668562, 0.00015502283, -9.377647e-06, -0.00038868943, 0.00014910729, -1.0255432e-05, -0.00031395876, 0.0001428222, -1.1014833e-05, -0.00024281604, 0.00013622786, -1.1660528e-05, -0.00017538297, 0.00012938173, -1.2197443e-05, -0.000111752735, 0.00012233843, -1.2630701e-05, -5.1991512e-05, 0.000115149596, -1.2965595e-05, 3.8598264e-06, 0.0001078639, -1.3207535e-05, 5.5784116e-05, 0.000100526966, -1.336202e-05, 0.00010378627, 9.318135e-05, -1.3434604e-05, 0.00014789162, 8.5866566e-05, -1.3430861e-05, 0.00018814433, 7.86191e-05, -1.3356356e-05, 0.00022460577, 7.147244e-05, -1.3216618e-05, 0.00025735295, 6.445709e-05, -1.3017114e-05, 0.000286477, 5.760067e-05, -1.2763224e-05, 0.00031208163, 5.092797e-05, -1.2460223e-05, 0.00033428168, 4.4461e-05, -1.2113258e-05, 0.00035320176, 3.8219114e-05, -1.1727332e-05, 0.0003689748, 3.2219068e-05, -1.130729e-05, 0.0003817409, 2.6475142e-05, -1.0857803e-05, 0.00039164576, 2.0999243e-05, -1.038336e-05, 0.00039884, 1.5801006e-05, -9.888251e-06, 0.00040347752, 1.0887914e-05, -9.376569e-06, 0.00040571476, 6.26541e-06, -8.852195e-06, 0.0004057096, 1.9370207e-06, -8.318794e-06, 0.00040362042, -2.0955258e-06, -7.7798195e-06, 0.00039960523, -5.8321793e-06, -7.2384996e-06, 0.00039382093, -9.274447e-06, -6.6978437e-06, 0.00038642244, -1.2425272e-05, -6.160641e-06, 0.00037756216, -1.5288915e-05, -5.629461e-06, 0.0003673893, -1.787084e-05, -5.106657e-06, 0.00035604928, -2.0177593e-05, -4.59437e-06, 0.0003436833, -2.2216695e-05, -4.0945292e-06, 0.0003304279, -2.399653e-05, -3.6088627e-06, 0.00031641452, -2.5526242e-05, -3.1388988e-06, 0.00030176924, -2.6815627e-05, -2.6859743e-06, 0.0002866125, -2.7875041e-05, -2.2512406e-06, 0.00027105885, -2.8715302e-05, -1.8356716e-06, 0.0002552167, -2.93476e-05, -1.4400705e-06, 0.00023918838, -2.9783418e-05, -1.0650791e-06, 0.00022306982, -3.0034436e-05, -7.1118507e-07, 0.00020695067, -3.0112476e-05, -3.7873096e-07, 0.00019091422, -3.0029418e-05, -6.792269e-08, 0.00017503738, -2.9797127e-05, 2.2116166e-07, 0.00015939082, -2.942741e-05, 4.885631e-07, 0.00014403896, -2.8931947e-05, 7.34433e-07, 0.00012904014, -2.832224e-05, 9.590243e-07, 0.00011444671, -2.7609563e-05, 1.162683e-06, 0.00010030521, -2.6804932e-05, 1.3458396e-06, 8.665654e-05, -2.5919051e-05, 1.5090006e-06, 7.353612e-05, -2.4962283e-05, 1.652741e-06, 6.0974133e-05, -2.3944629e-05, 1.7776961e-06, 4.8995713e-05, -2.2875689e-05, 1.8845531e-06, 3.762119e-05, -2.1764648e-05, 1.974045e-06, 2.6866323e-05, -2.0620257e-05, 2.0469433e-06, 1.6742535e-05, -1.9450816e-05, 2.1040503e-06, 7.2571747e-06, -1.8264162e-05, 2.1461933e-06, -1.5862436e-06, -1.706767e-05, 2.174219e-06, -9.787776e-06, -1.5868234e-05, 2.1889869e-06, -1.73508e-05, -1.467228e-05, 2.1913643e-06, -2.4281757e-05, -1.348575e-05, 2.182221e-06, -3.0589905e-05, -1.2314121e-05, 2.1624248e-06, -3.6287067e-05, -1.1162398e-05, 2.1328372e-06, -4.1387386e-05, -1.0035128e-05, 2.0943091e-06, -4.590709e-05, -8.936409e-06, 2.047677e-06, -4.9864255e-05, -7.869898e-06, 1.9937604e-06, -5.3278585e-05, -6.838821e-06, 1.9333577e-06, -5.6171193e-05, -5.8459955e-06, 1.8672445e-06, -5.856438e-05, -4.893837e-06, 1.7961705e-06, -6.048145e-05, -3.984378e-06, 1.7208582e-06, -6.194651e-05, -3.1192862e-06, 1.642e-06, -6.29843e-05, -2.2998786e-06, 1.5602578e-06, -6.3619984e-05, -1.5271424e-06, 1.4762613e-06, -6.3879044e-05, -8.017521e-07, 1.3906066e-06, -6.378706e-05, -1.2408844e-07, 1.3038565e-06, -6.336965e-05, 5.057424e-07, 1.2165387e-06, -6.2652245e-05, 1.0878899e-06, 1.129147e-06, -6.1660045e-05, 1.6227401e-06, 1.0421397e-06, -6.0417864e-05, 2.1108972e-06, 9.559409e-07, -5.8950045e-05, 2.553164e-06, 8.709398e-07, -5.728036e-05, 2.9505243e-06, 7.874921e-07, -5.5431923e-05, 3.3041247e-06, 7.059198e-07, -5.3427135e-05, 3.615257e-06, 6.265122e-07, -5.1287603e-05, 3.8853404e-06, 5.495268e-07, -4.9034094e-05, 4.1159074e-06, 4.751902e-07, -4.668647e-05, 4.3085847e-06, 4.0369903e-07, -4.4263674e-05, 4.46508e-06, 3.3522107e-07, -4.178368e-05, 4.5871666e-06, 2.6989662e-07, -3.9263476e-05, 4.67667e-06, 2.0783946e-07, -3.6719044e-05, 4.7354547e-06, 1.4913842e-07, -3.4165347e-05, 4.7654103e-06, 9.385847e-08, -3.161633e-05, 4.7684425e-06, 4.2042252e-08, -2.9084917e-05, 4.7464605e-06, -6.2886314e-09, -2.6583013e-05, 4.7013655e-06, -5.1132222e-08, -2.412152e-05, 4.635045e-06, -9.25048e-08, -2.1710353e-05, 4.5493603e-06, -1.3043949e-07, -1.9358455e-05, 4.446141e-06, -1.6498491e-07, -1.707382e-05, 4.327176e-06, -1.9620379e-07, -1.48635245e-05, 4.1942108e-06, -2.2417167e-07, -1.2733751e-05, 4.0489354e-06, -2.4897557e-07, -1.068982e-05, 3.8929857e-06, -2.707127e-07, -8.736229e-06, 3.7279349e-06, -2.8948926e-07, -6.8766813e-06, 3.5552912e-06, -3.0541926e-07, -5.1141283e-06, 3.376495e-06, -3.1862334e-07, -3.4508062e-06, 3.1929148e-06, -3.2922767e-07, -1.8882753e-06, 3.0058475e-06, -3.373629e-07, -4.2746012e-07, 2.8165139e-06, -3.431632e-07, 9.313091e-07, 2.6260607e-06, -3.467653e-07, 2.1882565e-06, 2.4355575e-06, -3.4830745e-07, 3.3441192e-06, 2.2459985e-06, -3.479289e-07, 4.4001076e-06, 2.0583013e-06, -3.4576885e-07, 5.3578647e-06, 1.8733089e-06, -3.419658e-07, 6.2194263e-06, 1.6917894e-06, -3.3665688e-07, 6.9871835e-06, 1.5144384e-06, -3.2997727e-07, 7.6638435e-06, 1.34188e-06, -3.2205966e-07, 8.252394e-06, 1.1746687e-06, -3.1303358e-07, 8.7560675e-06, 1.0132917e-06, -3.030252e-07, 9.178306e-06, 8.581711e-07, -2.921566e-07, 9.522731e-06, 7.0966644e-07, -2.8054586e-07, 9.793106e-06, 5.680768e-07, -2.6830622e-07, 9.993314e-06, 4.336444e-07, -2.555463e-07, 1.0127325e-05, 3.0655667e-07, -2.423695e-07, 1.0199168e-05, 1.8694958e-07, -2.2887416e-07, 1.0212908e-05, 7.4910524e-08, -2.1515312e-07, 1.0172623e-05, -2.95187e-08, -2.0129382e-07, 1.0082377e-05, -1.2633883e-07, -1.8737816e-07, 9.946208e-06, -2.1559009e-07, -1.734825e-07, 9.7680995e-06, -2.9734917e-07, -1.5967763e-07, 9.5519745e-06, -3.7172623e-07, -1.4602877e-07, 9.301667e-06, -4.3886186e-07, -1.3259574e-07, 9.02092e-06, -4.9892435e-07, -1.1943293e-07, 8.713363e-06, -5.5210666e-07, -1.0658943e-07, 8.38251e-06, -5.986237e-07, -9.41092e-08, 8.031741e-06, -6.3870976e-07, -8.203113e-08, 7.664302e-06, -6.726157e-07, -7.038927e-08, 7.2832904e-06, -7.006067e-07, -5.921297e-08, 6.8916556e-06, -7.229596e-07, -4.8527053e-08, 6.49219e-06, -7.399609e-07, -3.835203e-08, 6.087528e-06, -7.519044e-07, -2.8704285e-08, 5.680143e-06, -7.590891e-07, -1.9596296e-08, 5.2723453e-06, -7.618176e-07, -1.1036846e-08, 4.8662823e-06, -7.603939e-07, -3.031237e-09, 4.46394e-06, -7.551218e-07, 4.418483e-09, 4.067143e-06, -7.463035e-07, 1.1313302e-08, 3.677556e-06, -7.3423803e-07, 1.765702e-08, 3.2966882e-06, -7.1922e-07, 2.3456032e-08, 2.9258956e-06, -7.015382e-07, 2.8719102e-08, 2.5663846e-06, -6.814747e-07, 3.345716e-08, 2.2192173e-06, -6.5930385e-07, 3.7683073e-08, 1.8853157e-06, -6.3529126e-07, 4.1411457e-08, 1.565467e-06, -6.096932e-07, 4.4658474e-08, 1.2603292e-06, -5.827559e-07, 4.7441624e-08, 9.70437e-07, -5.5471486e-07, 4.9779572e-08, 6.9620745e-07, -5.2579463e-07, 5.169196e-08, 4.379468e-07, -4.962082e-07, 5.3199244e-08, 1.9585623e-07, -4.6615688e-07, 5.432252e-08, -2.9961402e-08, -4.3582997e-07, 5.5083376e-08, -2.3949508e-07, -4.054047e-07, 5.5503733e-08, -4.328192e-07, -3.7504617e-07, 5.5605728e-08, -6.1008706e-07, -3.449073e-07, 5.541156e-08, -7.715244e-07, -3.15129e-07, 5.4943396e-08, -9.174231e-07, -2.858402e-07, 5.422322e-08, -1.0481349e-06, -2.5715812e-07, 5.327278e-08, -1.1640653e-06, -2.2918846e-07, 5.2113457e-08, -1.2656678e-06, -2.020256e-07, 5.0766186e-08, -1.3534377e-06, -1.7575307e-07, 4.9251387e-08, -1.4279069e-06, -1.5044378e-07, 4.7588898e-08, -1.4896384e-06, -1.2616042e-07, 4.57979e-08, -1.5392213e-06, -1.0295587e-07, 4.3896875e-08, -1.5772656e-06, -8.087366e-08, 4.1903558e-08, -1.6043977e-06, -5.9948356e-08, 3.9834894e-08, -1.6212558e-06, -4.020604e-08, 3.770701e-08, -1.6284863e-06, -2.1664802e-08, 3.553519e-08, -1.6267392e-06, -4.335192e-09, 3.333386e-08, -1.6166646e-06, 1.1779286e-08, 3.1116556e-08, -1.5989098e-06, 2.6681693e-08, 2.8895943e-08, -1.5741152e-06, 4.0381167e-08, 2.6683795e-08, -1.5429129e-06, 5.2892442e-08, 2.4490996e-08, -1.5059222e-06, 6.423538e-08, 2.232756e-08, -1.463749e-06, 7.4434475e-08, 2.0202629e-08, -1.4169823e-06, 8.3518444e-08, 1.812449e-08, -1.3661931e-06, 9.151972e-08, 1.6100602e-08, -1.3119329e-06, 9.847406e-08, 1.4137604e-08, -1.2547313e-06, 1.044201e-07, 1.2241346e-08, -1.1950956e-06, 1.0939896e-07, 1.0416913e-08, -1.1335094e-06, 1.1345385e-07, 8.668654e-09, -1.0704321e-06, 1.1662968e-07, 7.0002133e-09, -1.0062978e-06, 1.1897273e-07, 5.4145577e-09, -9.415153e-07, 1.205303e-07, 3.914013e-09, -8.764674e-07, 1.2135041e-07, 2.5002977e-09, -8.1151114e-07, 1.2148145e-07, 1.1745553e-09, -7.469774e-07, 1.2097196e-07, -6.2609085e-11, -6.8317127e-07, 1.1987032e-07, -1.2110938e-09, -6.2037236e-07, 1.1822456e-07, -2.271265e-09, -5.58835e-07, 1.1608208e-07, -3.2439216e-09, -4.987888e-07, 1.13489484e-07, -4.13026e-09, -4.404392e-07, 1.1049239e-07, -4.9318403e-09, -3.839683e-07, 1.0713526e-07, -5.6505502e-09, -3.2953534e-07, 1.0346125e-07, -6.288575e-09, -2.772775e-07, 9.9512064e-08, -6.848361e-09, -2.27311e-07, 9.53279e-08, -7.332588e-09, -1.7973183e-07, 9.094725e-08, -7.744136e-09, -1.3461666e-07, 8.640693e-08, -8.086057e-09, -9.202395e-08, 8.1741916e-08, -8.361548e-09, -5.199485e-08, 7.698536e-08, -8.573921e-09, -1.45542485e-08, 7.2168504e-08, -8.726581e-09, 2.0288182e-08, 6.732069e-08, -8.822998e-09, 5.2536965e-08, 6.246931e-08, -8.86669e-09, 8.220977e-08, 5.763983e-08, -8.861194e-09, 1.09336405e-07, 5.2855775e-08, -8.81005e-09, 1.3395776e-07, 4.8138755e-08, -8.7167855e-09, 1.5612481e-07, 4.3508496e-08, -8.584893e-09, 1.7589768e-07, 3.898285e-08, -8.417816e-09, 1.9334462e-07, 3.457787e-08, -8.218936e-09, 2.0854107e-07, 3.0307817e-08, -7.991557e-09, 2.2156881e-07, 2.618524e-08, -7.738895e-09, 2.3251502e-07, 2.2221032e-08, -7.464069e-09, 2.414715e-07, 1.8424474e-08, -7.17009e-09, 2.4853378e-07, 1.4803324e-08, -6.8598527e-09, 2.538005e-07, 1.13638645e-08, -6.5361303e-09, 2.5737245e-07, 8.110991e-09, -6.201568e-09, 2.5935213e-07, 5.04828e-09, -5.8586775e-09, 2.59843e-07, 2.1780626e-09, -5.509836e-09, 2.589488e-07, -4.9849536e-10, -5.15728e-09, 2.567731e-07, -2.981318e-09, -4.8031072e-09, 2.534187e-07, -5.271341e-09, -4.4492725e-09, 2.4898725e-07, -7.3704363e-09, -4.0975907e-09, 2.4357865e-07, -9.281332e-09, -3.749735e-09, 2.372908e-07, -1.1007541e-08, -3.4072398e-09, 2.3021916e-07, -1.2553282e-08, -3.0715013e-09, 2.2245644e-07, -1.3923415e-08, -2.7437814e-09, 2.1409232e-07, -1.5123362e-08, -2.4252103e-09, 2.0521321e-07, -1.615904e-08, -2.1167894e-09, 1.9590203e-07, -1.7036802e-08, -1.8193966e-09, 1.86238e-07, -1.7763364e-08, -1.5337895e-09, 1.7629652e-07, -1.834575e-08, -1.2606101e-09, 1.6614908e-07, -1.8791228e-08, -1.0003902e-09, 1.5586309e-07, -1.9107263e-08, -7.5355633e-10, 1.4550189e-07, -1.9301458e-08, -5.20435e-10, 1.3512468e-07, -1.9381504e-08, -3.01258e-10, 1.2478652e-07, -1.9355136e-08, -9.616834e-11, 1.1453834e-07, -1.9230091e-08, 9.477451e-11, 1.04426945e-07, -1.9014069e-08, 2.7158878e-10, 9.4495114e-08, -1.8714683e-08, 4.3436485e-10, 8.478162e-08, -1.8339447e-08, 5.8325955e-10, 7.5321324e-08, -1.7895728e-08, 7.184906e-10, 6.614531e-08, -1.7390718e-08, 8.403312e-10, 5.728095e-08, -1.683142e-08, 9.491047e-10, 4.8752035e-08, -1.6224616e-08, 1.0451789e-09, 4.0578925e-08, -1.5576854e-08, 1.1289618e-09, 3.2778672e-08, -1.4894421e-08, 1.2008959e-09, 2.5365173e-08, -1.418334e-08, 1.2614535e-09, 1.8349327e-08, -1.3449352e-08, 1.3111325e-09, 1.1739186e-08, -1.2697905e-08, 1.3504518e-09, 5.5401195e-09, -1.19341514e-08, 1.3799466e-09, -2.4502214e-10, -1.1162937e-08, 1.4001657e-09, -5.615743e-09, -1.0388803e-08, 1.4116661e-09, -1.0573735e-08, -9.615977e-09, 1.415011e-09, -1.5122714e-08, -8.848384e-09, 1.4107654e-09, -1.9268256e-08, -8.0896365e-09, 1.3994932e-09, -2.3017634e-08, -7.3430453e-09, 1.381755e-09, -2.6379661e-08, -6.6116215e-09, 1.3581047e-09, -2.936453e-08, -5.8980816e-09, 1.3290873e-09, -3.198367e-08, -5.2048557e-09, 1.2952369e-09, -3.424959e-08, -4.534095e-09, 1.2570746e-09, -3.617575e-08, -3.8876795e-09, 1.2151063e-09, -3.7776395e-08, -3.2672298e-09, 1.1698224e-09, -3.9066464e-08, -2.6741145e-09, 1.1216944e-09, -4.006143e-08, -2.1094635e-09, 1.0711757e-09, -4.0777202e-08, -1.5741773e-09, 1.0186996e-09, -4.1229995e-08, -1.0689402e-09, 9.646783e-10, -4.143624e-08, -5.942309e-10, 9.095031e-10, -4.1412477e-08, -1.503358e-10, 8.5354285e-10, -4.1175248e-08, 2.626395e-10, 7.971444e-10, -4.0741035e-08, 6.4475747e-10, 7.4063206e-10, -4.012616e-08, 9.962365e-10, 6.843076e-10, -3.934672e-08, 1.3174387e-09, 6.284503e-10, -3.841852e-08, 1.6088574e-09, 5.733169e-10, -3.7357e-08, 1.8711055e-09, 5.191422e-10, -3.6177198e-08, 2.1049036e-09, 4.661391e-10, -3.4893695e-08, 2.311069e-09, 4.1449952e-10, -3.3520564e-08, 2.4905038e-09, 3.6439418e-10, -3.2071334e-08, 2.6441846e-09, 3.1597394e-10, -3.055898e-08, 2.7731526e-09, 2.6936997e-10, -2.8995856e-08, 2.878502e-09, 2.2469474e-10, -2.7393716e-08, 2.961373e-09, 1.8204259e-10, -2.5763667e-08, 3.0229395e-09, 1.4149064e-10, -2.4116174e-08, 3.0644036e-09, 1.03099605e-10, -2.2461041e-08, 3.0869853e-09, 6.691461e-11, -2.0807413e-08, 3.091916e-09, 3.2966126e-11, -1.9163773e-08, 3.0804304e-09, 1.2708049e-12, -1.7537948e-08, 3.0537604e-09, -2.8167592e-11, -1.5937113e-08, 3.0131293e-09, -5.5357295e-11, -1.43678e-08, 2.9597451e-09, -8.031763e-11, -1.2835912e-08, 2.894796e-09, -1.0307812e-10, -1.1346734e-08, 2.8194451e-09, -1.2367762e-10, -9.904955e-09, 2.734827e-09, -1.4216345e-10, -8.514679e-09, 2.6420433e-09, -1.5859047e-10, -7.1794513e-09, 2.5421587e-09, -1.7302042e-10, -5.9022778e-09, 2.4361997e-09, -1.855209e-10, -4.685649e-09, 2.3251503e-09, -1.9616479e-10, -3.5315615e-09, 2.209951e-09, -2.0502935e-10, -2.4415447e-09, 2.0914972e-09, -2.1219564e-10, -1.4166869e-09, 1.9706363e-09, -2.1774765e-10, -4.5765883e-10, 1.8481682e-09, -2.2177188e-10, 4.3525783e-10, 1.7248439e-09, -2.2435648e-10, 1.2621453e-09, 1.6013654e-09, -2.2559085e-10, 2.023423e-09, 1.4783852e-09, -2.2556501e-10, 2.7198213e-09, 1.3565067e-09, -2.2436909e-10, 3.3523553e-09, 1.2362844e-09, -2.2209286e-10, 3.9222994e-09, 1.1182247e-09, -2.188253e-10, 4.4311625e-09, 1.0027865e-09, -2.1465418e-10, 4.880663e-09, 8.9038227e-10, -2.0966572e-10, 5.272705e-09, 7.8137946e-10, -2.0394417e-10, 5.6093548e-09, 6.761014e-10, -1.9757164e-10, 5.892819e-09, 5.7482913e-10, -1.9062771e-10, 6.1254233e-09, 4.778027e-10, -1.8318927e-10};
	localparam real hb[0:1199] = {0.024535134, 0.00031300698, -0.0002562084, 0.024466371, 0.00044678675, -0.00025098654, 0.024331018, 0.000577397, -0.00024344047, 0.024130605, 0.00070377014, -0.00023387383, 0.023867166, 0.0008249804, -0.0002225721, 0.023543173, 0.00094023533, -0.00020980298, 0.023161484, 0.0010488675, -0.00019581664, 0.022725265, 0.0011503266, -0.0001808461, 0.022237957, 0.0012441713, -0.00016510769, 0.021703204, 0.0013300614, -0.00014880144, 0.021124823, 0.0014077503, -0.00013211157, 0.020506745, 0.0014770778, -0.000115206974, 0.019852985, 0.0015379628, -9.824172e-05, 0.019167598, 0.0015903963, -8.135559e-05, 0.01845465, 0.0016344344, -6.467463e-05, 0.017718183, 0.001670193, -4.831171e-05, 0.016962186, 0.0016978399, -3.236711e-05, 0.016190572, 0.0017175906, -1.6929074e-05, 0.015407158, 0.0017297013, -2.0744324e-06, 0.014615638, 0.0017344642, 1.21308285e-05, 0.013819575, 0.0017322025, 2.5630961e-05, 0.013022378, 0.0017232649, 3.837986e-05, 0.012227292, 0.0017080221, 5.034048e-05, 0.011437392, 0.0016868612, 6.148425e-05, 0.010655567, 0.001660183, 7.179047e-05, 0.009884519, 0.0016283974, 8.1245795e-05, 0.0091267545, 0.0015919203, 8.984361e-05, 0.008384588, 0.0015511703, 9.7583536e-05, 0.00766013, 0.0015065657, 0.00010447088, 0.0069552967, 0.0014585223, 0.000110516085, 0.006271805, 0.0014074501, 0.000115734285, 0.005611177, 0.0013537516, 0.000120144796, 0.004974743, 0.0012978201, 0.00012377062, 0.0043636453, 0.0012400375, 0.00012663804, 0.0037788455, 0.0011807726, 0.00012877617, 0.0032211267, 0.0011203804, 0.00013021656, 0.0026911027, 0.0010592001, 0.00013099279, 0.0021892241, 0.0009975553, 0.0001311401, 0.0017157864, 0.00093575194, 0.00013069507, 0.0012709373, 0.00087407854, 0.0001296953, 0.0008546855, 0.00081280543, 0.00012817905, 0.0004669088, 0.00075218437, 0.000126185, 0.00010736289, 0.00069244846, 0.00012375199, -0.00022430973, 0.00063381204, 0.00012091877, -0.0005285711, 0.00057647086, 0.000117723765, -0.00080597884, 0.0005206019, 0.00011420487, -0.0010571777, 0.00046636406, 0.0001103993, -0.0012828903, 0.00041389815, 0.000106343374, -0.0014839094, 0.0003633275, 0.000102072416, -0.0016610889, 0.0003147584, 9.7620585e-05, -0.0018153363, 0.00026828056, 9.302079e-05, -0.0019476044, 0.00022396795, 8.830458e-05, -0.002058884, 0.00018187916, 8.350206e-05, -0.0021501961, 0.00014205833, 7.864182e-05, -0.0022225862, 0.00010453572, 7.375089e-05, -0.0022771163, 6.9328555e-05, 6.88547e-05, -0.0023148593, 3.644175e-05, 6.3977044e-05, -0.0023368932, 5.8687147e-06, 5.914005e-05, -0.002344295, -2.2407867e-05, 5.4364198e-05, -0.0023381358, -4.841523e-05, 4.966832e-05, -0.0023194766, -7.2189745e-05, 4.5069588e-05, -0.0022893632, -9.377611e-05, 4.0583553e-05, -0.0022488215, -0.00011322658, 3.6224174e-05, -0.0021988559, -0.00013060021, 3.200384e-05, -0.0021404433, -0.00014596208, 2.7933427e-05, -0.0020745327, -0.0001593826, 2.4022327e-05, -0.0020020404, -0.00017093674, 2.0278512e-05, -0.0019238496, -0.00018070341, 1.6708584e-05, -0.0018408066, -0.00018876477, 1.3317829e-05, -0.0017537207, -0.00019520559, 1.0110291e-05, -0.001663362, -0.00020011268, 7.088825e-06, -0.0015704606, -0.00020357428, 4.255167e-06, -0.0014757058, -0.00020567955, 1.61e-06, -0.0013797453, -0.00020651803, -8.4697547e-07, -0.0012831856, -0.00020617925, -3.1169748e-06, -0.0011865911, -0.00020475216, -5.2020596e-06, -0.0010904848, -0.00020232481, -7.1050695e-06, -0.0009953484, -0.00019898398, -8.829555e-06, -0.0009016233, -0.00019481475, -1.0379707e-05, -0.0008097103, -0.00018990033, -1.17602995e-05, -0.00071997166, -0.00018432162, -1.2976615e-05, -0.0006327311, -0.00017815706, -1.4034391e-05, -0.00054827565, -0.0001714824, -1.4939754e-05, -0.0004668562, -0.00016437052, -1.5699165e-05, -0.00038868943, -0.00015689118, -1.631936e-05, -0.00031395876, -0.00014911102, -1.6807302e-05, -0.00024281604, -0.00014109333, -1.7170125e-05, -0.00017538297, -0.00013289804, -1.7415086e-05, -0.000111752735, -0.00012458164, -1.7549526e-05, -5.1991512e-05, -0.00011619707, -1.7580818e-05, 3.8598264e-06, -0.000107793836, -1.7516333e-05, 5.5784116e-05, -9.94179e-05, -1.7363402e-05, 0.00010378627, -9.111173e-05, -1.712928e-05, 0.00014789162, -8.291434e-05, -1.6821115e-05, 0.00018814433, -7.4861324e-05, -1.6445923e-05, 0.00022460577, -6.698494e-05, -1.6010556e-05, 0.00025735295, -5.931417e-05, -1.552168e-05, 0.000286477, -5.187481e-05, -1.4985756e-05, 0.00031208163, -4.468957e-05, -1.4409022e-05, 0.00033428168, -3.7778165e-05, -1.3797476e-05, 0.00035320176, -3.1157462e-05, -1.315686e-05, 0.0003689748, -2.4841554e-05, -1.2492656e-05, 0.0003817409, -1.8841929e-05, -1.1810067e-05, 0.00039164576, -1.3167571e-05, -1.1114017e-05, 0.00039884, -7.825109e-06, -1.0409144e-05, 0.00040347752, -2.8189438e-06, -9.6997965e-06, 0.00040571476, 1.8486062e-06, -8.9900295e-06, 0.0004057096, 6.177173e-06, -8.28361e-06, 0.00040362042, 1.0168196e-05, -7.584015e-06, 0.00039960523, 1.3824786e-05, -6.8944314e-06, 0.00039382093, 1.7151588e-05, -6.2177664e-06, 0.00038642244, 2.0154645e-05, -5.556649e-06, 0.00037756216, 2.2841263e-05, -4.913437e-06, 0.0003673893, 2.5219893e-05, -4.2902248e-06, 0.00035604928, 2.729999e-05, -3.6888503e-06, 0.0003436833, 2.90919e-05, -3.1109055e-06, 0.0003304279, 3.0606734e-05, -2.5577447e-06, 0.00031641452, 3.185627e-05, -2.0304954e-06, 0.00030176924, 3.285283e-05, -1.5300673e-06, 0.0002866125, 3.360917e-05, -1.0571654e-06, 0.00027105885, 3.4138407e-05, -6.122993e-07, 0.0002552167, 3.4453897e-05, -1.9579534e-07, 0.00023918838, 3.4569166e-05, 1.9219195e-07, 0.00022306982, 3.4497825e-05, 5.516684e-07, 0.00020695067, 3.425348e-05, 8.827886e-07, 0.00019091422, 3.384968e-05, 1.1858444e-06, 0.00017503738, 3.329983e-05, 1.4612535e-06, 0.00015939082, 3.2617154e-05, 1.7095485e-06, 0.00014403896, 3.1814616e-05, 1.9313652e-06, 0.00012904014, 3.090489e-05, 2.1274325e-06, 0.00011444671, 2.9900291e-05, 2.2985619e-06, 0.00010030521, 2.8812772e-05, 2.4456365e-06, 8.665654e-05, 2.7653854e-05, 2.5696029e-06, 7.353612e-05, 2.6434613e-05, 2.67146e-06, 6.0974133e-05, 2.516565e-05, 2.7522506e-06, 4.8995713e-05, 2.3857068e-05, 2.8130535e-06, 3.762119e-05, 2.2518461e-05, 2.8549744e-06, 2.6866323e-05, 2.1158894e-05, 2.8791387e-06, 1.6742535e-05, 1.9786898e-05, 2.886684e-06, 7.2571747e-06, 1.841046e-05, 2.878753e-06, -1.5862436e-06, 1.7037019e-05, 2.8564882e-06, -9.787776e-06, 1.5673473e-05, 2.821025e-06, -1.73508e-05, 1.4326178e-05, 2.7734864e-06, -2.4281757e-05, 1.3000951e-05, 2.714978e-06, -3.0589905e-05, 1.1703081e-05, 2.6465846e-06, -3.6287067e-05, 1.0437339e-05, 2.5693641e-06, -4.1387386e-05, 9.20799e-06, 2.4843455e-06, -4.590709e-05, 8.018806e-06, 2.3925247e-06, -4.9864255e-05, 6.873081e-06, 2.2948623e-06, -5.3278585e-05, 5.7736515e-06, 2.1922804e-06, -5.6171193e-05, 4.7229096e-06, 2.0856617e-06, -5.856438e-05, 3.7228258e-06, 1.975846e-06, -6.048145e-05, 2.7749675e-06, 1.8636309e-06, -6.194651e-05, 1.8805188e-06, 1.7497688e-06, -6.29843e-05, 1.0403033e-06, 1.6349672e-06, -6.3619984e-05, 2.5480426e-07, 1.5198887e-06, -6.3879044e-05, -4.7581312e-07, 1.4051493e-06, -6.378706e-05, -1.15168e-06, 1.2913197e-06, -6.336965e-05, -1.773202e-06, 1.1789253e-06, -6.2652245e-05, -2.3410378e-06, 1.0684464e-06, -6.1660045e-05, -2.8560773e-06, 9.603193e-07, -6.0417864e-05, -3.319421e-06, 8.549368e-07, -5.8950045e-05, -3.7323584e-06, 7.5264956e-07, -5.728036e-05, -4.096349e-06, 6.537673e-07, -5.5431923e-05, -4.4130024e-06, 5.585597e-07, -5.3427135e-05, -4.6840573e-06, 4.6725842e-07, -5.1287603e-05, -4.9113664e-06, 3.8005817e-07, -4.9034094e-05, -5.0968765e-06, 2.971185e-07, -4.668647e-05, -5.242612e-06, 2.1856553e-07, -4.4263674e-05, -5.35066e-06, 1.4449361e-07, -4.178368e-05, -5.423153e-06, 7.496708e-08, -3.9263476e-05, -5.462257e-06, 1.002211e-08, -3.6719044e-05, -5.470155e-06, -5.033148e-08, -3.4165347e-05, -5.4490374e-06, -1.06108395e-07, -3.161633e-05, -5.4010884e-06, -1.5734604e-07, -2.9084917e-05, -5.3284753e-06, -2.0410272e-07, -2.6583013e-05, -5.233338e-06, -2.464558e-07, -2.412152e-05, -5.117782e-06, -2.8450006e-07, -2.1710353e-05, -4.9838673e-06, -3.1834574e-07, -1.9358455e-05, -4.833602e-06, -3.4811717e-07, -1.707382e-05, -4.668936e-06, -3.7395077e-07, -1.48635245e-05, -4.491755e-06, -3.9599382e-07, -1.2733751e-05, -4.303874e-06, -4.1440268e-07, -1.068982e-05, -4.107035e-06, -4.2934144e-07, -8.736229e-06, -3.9029005e-06, -4.4098041e-07, -6.8766813e-06, -3.6930542e-06, -4.4949502e-07, -5.1141283e-06, -3.4789944e-06, -4.5506425e-07, -3.4508062e-06, -3.2621354e-06, -4.5786967e-07, -1.8882753e-06, -3.0438046e-06, -4.5809418e-07, -4.2746012e-07, -2.825242e-06, -4.5592108e-07, 9.313091e-07, -2.6076007e-06, -4.51533e-07, 2.1882565e-06, -2.3919458e-06, -4.45111e-07, 3.3441192e-06, -2.1792569e-06, -4.3683377e-07, 4.4001076e-06, -1.9704275e-06, -4.2687697e-07, 5.3578647e-06, -1.7662677e-06, -4.1541227e-07, 6.2194263e-06, -1.567505e-06, -4.0260707e-07, 6.9871835e-06, -1.3747872e-06, -3.8862368e-07, 7.6638435e-06, -1.1886843e-06, -3.7361895e-07, 8.252394e-06, -1.0096911e-06, -3.5774383e-07, 8.7560675e-06, -8.3823016e-07, -3.4114302e-07, 9.178306e-06, -6.7465476e-07, -3.2395465e-07, 9.522731e-06, -5.1925196e-07, -3.0631003e-07, 9.793106e-06, -3.7224575e-07, -2.883335e-07, 9.993314e-06, -2.3380052e-07, -2.7014212e-07, 1.0127325e-05, -1.0402444e-07, -2.5184588e-07, 1.0199168e-05, 1.7027123e-08, -2.335473e-07, 1.0212908e-05, 1.293481e-07, -2.1534167e-07, 1.0172623e-05, 2.329782e-07, -1.9731698e-07, 1.0082377e-05, 3.2799952e-07, -1.7955396e-07, 9.946208e-06, 4.1453296e-07, -1.6212627e-07, 9.7680995e-06, 4.92735e-07, -1.4510051e-07, 9.5519745e-06, 5.627941e-07, -1.2853647e-07, 9.301667e-06, 6.249278e-07, -1.1248726e-07, 9.02092e-06, 6.7937896e-07, -9.699951e-08, 8.713363e-06, 7.2641336e-07, -8.21136e-08, 8.38251e-06, 7.6631613e-07, -6.7863915e-08, 8.031741e-06, 7.9938917e-07, -5.427908e-08, 7.664302e-06, 8.259483e-07, -4.1382197e-08, 7.2832904e-06, 8.4632063e-07, -2.919116e-08, 6.8916556e-06, 8.608421e-07, -1.7718913e-08, 6.49219e-06, 8.6985494e-07, -6.97374e-09, 6.087528e-06, 8.737057e-07, 3.0404461e-09, 5.680143e-06, 8.72743e-07, 1.2323809e-08, 5.2723453e-06, 8.673155e-07, 2.0880298e-08, 4.8662823e-06, 8.577702e-07, 2.871736e-08, 4.46394e-06, 8.444507e-07, 3.5845645e-08, 4.067143e-06, 8.276957e-07, 4.2278728e-08, 3.677556e-06, 8.078376e-07, 4.803283e-08, 3.2966882e-06, 7.8520105e-07, 5.3126534e-08, 2.9258956e-06, 7.6010207e-07, 5.7580532e-08, 2.5663846e-06, 7.328469e-07, 6.141737e-08, 2.2192173e-06, 7.0373113e-07, 6.4661165e-08, 1.8853157e-06, 6.730388e-07, 6.7337425e-08, 1.565467e-06, 6.41042e-07, 6.9472776e-08, 1.2603292e-06, 6.0800005e-07, 7.109473e-08, 9.70437e-07, 5.7415923e-07, 7.2231536e-08, 6.9620745e-07, 5.397524e-07, 7.291193e-08, 4.379468e-07, 5.049988e-07, 7.316496e-08, 1.9585623e-07, 4.7010366e-07, 7.3019834e-08, -2.9961402e-08, 4.3525836e-07, 7.2505735e-08, -2.3949508e-07, 4.0064037e-07, 7.1651684e-08, -4.328192e-07, 3.6641333e-07, 7.0486394e-08, -6.1008706e-07, 3.327271e-07, 6.903814e-08, -7.715244e-07, 2.9971807e-07, 6.733465e-08, -9.174231e-07, 2.675094e-07, 6.540301e-08, -1.0481349e-06, 2.3621119e-07, 6.326954e-08, -1.1640653e-06, 2.0592107e-07, 6.0959735e-08, -1.2656678e-06, 1.767244e-07, 5.849819e-08, -1.3534377e-06, 1.4869475e-07, 5.5908533e-08, -1.4279069e-06, 1.2189444e-07, 5.321336e-08, -1.4896384e-06, 9.6374876e-08, 5.043421e-08, -1.5392213e-06, 7.217718e-08, 4.7591517e-08, -1.5772656e-06, 4.9332662e-08, 4.4704592e-08, -1.6043977e-06, 2.7863374e-08, 4.1791584e-08, -1.6212558e-06, 7.782636e-09, 3.8869494e-08, -1.6284863e-06, -1.0904391e-08, 3.595415e-08, -1.6267392e-06, -2.8200155e-08, 3.306022e-08, -1.6166646e-06, -4.411416e-08, 3.0201203e-08, -1.5989098e-06, -5.8662405e-08, 2.7389465e-08, -1.5741152e-06, -7.186684e-08, 2.4636233e-08, -1.5429129e-06, -8.375485e-08, 2.1951633e-08, -1.5059222e-06, -9.435867e-08, 1.9344714e-08, -1.463749e-06, -1.03714925e-07, 1.6823469e-08, -1.4169823e-06, -1.1186411e-07, 1.439488e-08, -1.3661931e-06, -1.1885009e-07, 1.2064946e-08, -1.3119329e-06, -1.2471963e-07, 9.838728e-09, -1.2547313e-06, -1.29522e-07, 7.7203826e-09, -1.1950956e-06, -1.3330842e-07, 5.7132135e-09, -1.1335094e-06, -1.361318e-07, 3.8197085e-09, -1.0704321e-06, -1.3804626e-07, 2.0415873e-09, -1.0062978e-06, -1.3910675e-07, 3.7984801e-10, -9.415153e-07, -1.3936874e-07, -1.1651876e-09, -8.764674e-07, -1.388879e-07, -2.593827e-09, -8.1151114e-07, -1.377198e-07, -3.90696e-09, -7.469774e-07, -1.3591956e-07, -5.1060143e-09, -6.8317127e-07, -1.335417e-07, -6.192906e-09, -6.2037236e-07, -1.3063982e-07, -7.1699997e-09, -5.58835e-07, -1.2726642e-07, -8.040059e-09, -4.987888e-07, -1.234727e-07, -8.806209e-09, -4.404392e-07, -1.193084e-07, -9.471889e-09, -3.839683e-07, -1.1482161e-07, -1.0040816e-08, -3.2953534e-07, -1.1005868e-07, -1.0516945e-08, -2.772775e-07, -1.0506407e-07, -1.0904428e-08, -2.27311e-07, -9.9880275e-08, -1.1207582e-08, -1.7973183e-07, -9.4547744e-08, -1.1430856e-08, -1.3461666e-07, -8.91048e-08, -1.1578795e-08, -9.202395e-08, -8.358762e-08, -1.16560095e-08, -5.199485e-08, -7.803016e-08, -1.1667149e-08, -1.45542485e-08, -7.246417e-08, -1.16168755e-08, 2.0288182e-08, -6.6919185e-08, -1.1509836e-08, 5.2536965e-08, -6.1422504e-08, -1.13506395e-08, 8.220977e-08, -5.5999248e-08, -1.1143839e-08, 1.09336405e-07, -5.067234e-08, -1.0893908e-08, 1.3395776e-07, -4.5462585e-08, -1.0605226e-08, 1.5612481e-07, -4.0388677e-08, -1.028206e-08, 1.7589768e-07, -3.5467277e-08, -9.928551e-09, 1.9334462e-07, -3.0713068e-08, -9.548704e-09, 2.0854107e-07, -2.6138807e-08, -9.1463725e-09, 2.2156881e-07, -2.175541e-08, -8.725253e-09, 2.3251502e-07, -1.757202e-08, -8.288875e-09, 2.414715e-07, -1.3596089e-08, -7.840597e-09, 2.4853378e-07, -9.8334585e-09, -7.3835946e-09, 2.538005e-07, -6.288444e-09, -6.920868e-09, 2.5737245e-07, -2.9639238e-09, -6.4552292e-09, 2.5935213e-07, 1.385764e-10, -5.989305e-09, 2.59843e-07, 3.018793e-09, -5.5255374e-09, 2.589488e-07, 5.677636e-09, -5.0661817e-09, 2.567731e-07, 8.117101e-09, -4.613309e-09, 2.534187e-07, 1.034018e-08, -4.1688093e-09, 2.4898725e-07, 1.2350776e-08, -3.7343946e-09, 2.4357865e-07, 1.4153619e-08, -3.3116012e-09, 2.372908e-07, 1.5754177e-08, -2.9017961e-09, 2.3021916e-07, 1.715858e-08, -2.5061806e-09, 2.2245644e-07, 1.8373541e-08, -2.125797e-09, 2.1409232e-07, 1.9406276e-08, -1.761534e-09, 2.0521321e-07, 2.0264434e-08, -1.4141326e-09, 1.9590203e-07, 2.0956023e-08, -1.0841935e-09, 1.86238e-07, 2.1489345e-08, -7.721841e-10, 1.7629652e-07, 2.1872934e-08, -4.7844484e-10, 1.6614908e-07, 2.2115486e-08, -2.0319714e-10, 1.5586309e-07, 2.2225818e-08, 5.344951e-11, 1.4550189e-07, 2.2212795e-08, 2.9149008e-10, 1.3512468e-07, 2.2085295e-08, 5.110166e-10, 1.2478652e-07, 2.1852157e-08, 7.122107e-10, 1.1453834e-07, 2.1522137e-08, 8.9533625e-10, 1.04426945e-07, 2.1103865e-08, 1.0607322e-09, 9.4495114e-08, 2.0605821e-08, 1.2088054e-09, 8.478162e-08, 2.0036286e-08, 1.3400235e-09, 7.5321324e-08, 1.9403327e-08, 1.4549087e-09, 6.614531e-08, 1.871476e-08, 1.5540305e-09, 5.728095e-08, 1.7978135e-08, 1.6379994e-09, 4.8752035e-08, 1.720071e-08, 1.7074615e-09, 4.0578925e-08, 1.6389441e-08, 1.7630918e-09, 3.2778672e-08, 1.5550954e-08, 1.8055891e-09, 2.5365173e-08, 1.46915555e-08, 1.8356706e-09, 1.8349327e-08, 1.3817201e-08, 1.8540666e-09, 1.1739186e-08, 1.29335e-08, 1.8615159e-09, 5.5401195e-09, 1.2045713e-08, 1.8587619e-09, -2.4502214e-10, 1.1158744e-08, 1.8465472e-09, -5.615743e-09, 1.0277143e-08, 1.8256112e-09, -1.0573735e-08, 9.405107e-09, 1.7966854e-09, -1.5122714e-08, 8.546483e-09, 1.7604905e-09, -1.9268256e-08, 7.704774e-09, 1.717734e-09, -2.3017634e-08, 6.883146e-09, 1.6691063e-09, -2.6379661e-08, 6.0844334e-09, 1.6152796e-09, -2.936453e-08, 5.3111493e-09, 1.5569047e-09, -3.198367e-08, 4.5654955e-09, 1.4946098e-09, -3.424959e-08, 3.849373e-09, 1.4289985e-09, -3.617575e-08, 3.1643923e-09, 1.3606484e-09, -3.7776395e-08, 2.5118894e-09, 1.2901102e-09, -3.9066464e-08, 1.8929347e-09, 1.2179068e-09, -4.006143e-08, 1.308348e-09, 1.1445321e-09, -4.0777202e-08, 7.587121e-10, 1.0704512e-09, -4.1229995e-08, 2.4438676e-10, 9.960991e-10, -4.143624e-08, -2.344776e-10, 9.218817e-10, -4.1412477e-08, -6.7792555e-10, 8.4817486e-10, -4.1175248e-08, -1.0861823e-09, 7.7532514e-10, -4.0741035e-08, -1.4596401e-09, 7.0364975e-10, -4.012616e-08, -1.7988436e-09, 6.334373e-10, -3.934672e-08, -2.1044768e-09, 5.6494803e-10, -3.841852e-08, -2.3773494e-09, 4.9841475e-10, -3.7357e-08, -2.6183833e-09, 4.3404344e-10, -3.6177198e-08, -2.8285996e-09, 3.7201414e-10, -3.4893695e-08, -3.0091072e-09, 3.1248187e-10, -3.3520564e-08, -3.16109e-09, 2.5557761e-10, -3.2071334e-08, -3.2857954e-09, 2.0140933e-10, -3.055898e-08, -3.3845236e-09, 1.5006307e-10, -2.8995856e-08, -3.4586167e-09, 1.01604045e-10, -2.7393716e-08, -3.509449e-09, 5.607785e-11, -2.5763667e-08, -3.5384178e-09, 1.3511569e-11, -2.4116174e-08, -3.5469339e-09, -2.6085033e-11, -2.2461041e-08, -3.5364134e-09, -6.271831e-11, -2.0807413e-08, -3.5082708e-09, -9.6409554e-11, -1.9163773e-08, -3.463911e-09, -1.2719384e-10, -1.7537948e-08, -3.404722e-09, -1.5511882e-10, -1.5937113e-08, -3.3320708e-09, -1.802436e-10, -1.43678e-08, -3.2472962e-09, -2.0263764e-10, -1.2835912e-08, -3.1517042e-09, -2.2237959e-10, -1.1346734e-08, -3.0465643e-09, -2.395563e-10, -9.904955e-09, -2.9331046e-09, -2.542617e-10, -8.514679e-09, -2.8125087e-09, -2.6659588e-10, -7.1794513e-09, -2.6859126e-09, -2.766641e-10, -5.9022778e-09, -2.5544027e-09, -2.8457592e-10, -4.685649e-09, -2.419013e-09, -2.9044417e-10, -3.5315615e-09, -2.2807243e-09, -2.9438432e-10, -2.4415447e-09, -2.140462e-09, -2.9651362e-10, -1.4166869e-09, -1.9990956e-09, -2.9695033e-10, -4.5765883e-10, -1.8574386e-09, -2.95813e-10, 4.3525783e-10, -1.7162478e-09, -2.9322003e-10, 1.2621453e-09, -1.5762234e-09, -2.892888e-10, 2.023423e-09, -1.4380094e-09, -2.8413527e-10, 2.7198213e-09, -1.3021949e-09, -2.7787359e-10, 3.3523553e-09, -1.169314e-09, -2.706154e-10, 3.9222994e-09, -1.0398475e-09, -2.6246955e-10, 4.4311625e-09, -9.142245e-10, -2.5354177e-10, 4.880663e-09, -7.928229e-10, -2.439343e-10, 5.272705e-09, -6.7597217e-10, -2.3374555e-10, 5.6093548e-09, -5.6395427e-10, -2.2307003e-10, 5.892819e-09, -4.5700616e-10, -2.1199795e-10, 6.1254233e-09, -3.5532136e-10, -2.0061512e-10};
endpackage
`endif
