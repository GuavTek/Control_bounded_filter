`ifndef COEFFICIENTS_FX_SV_
`define COEFFICIENTS_FX_SV_
package Coefficients_Fx;
	localparam N = 2;
	localparam M = 2;
	localparam COEFF_BIAS = 48;
	localparam logic signed[63:0] Lfr[0:1] = {64'd261916578309020, 64'd261916578309020};
	localparam logic signed[63:0] Lfi[0:1] = {64'd24304793653278, - 64'd24304793653278};
	localparam logic signed[63:0] Lbr[0:1] = {64'd261916578309020, 64'd261916578309020};
	localparam logic signed[63:0] Lbi[0:1] = {64'd24304793653278, - 64'd24304793653278};
	localparam logic signed[63:0] Wfr[0:1] = {- 64'd3161610580726, - 64'd3161610580726};
	localparam logic signed[63:0] Wfi[0:1] = {- 64'd4798877033583, 64'd4798877033583};
	localparam logic signed[63:0] Wbr[0:1] = {- 64'd3161610580726, - 64'd3161610580726};
	localparam logic signed[63:0] Wbi[0:1] = {- 64'd4798877033583, 64'd4798877033583};
	localparam logic signed[63:0] Ffr[0:1][0:39] = '{
		'{- 64'd16661173520135, - 64'd67604904587707, - 64'd46932306946327, - 64'd58666327761395, - 64'd72791968326060, - 64'd50139480307340, - 64'd94481366958141, - 64'd42076947065871, - 64'd112262382465842, - 64'd34518947358519, - 64'd126411729164527, - 64'd27494407471536, - 64'd137215677493413, - 64'd21022035995946, - 64'd144965326781880, - 64'd15111388452564, - 64'd149952417573864, - 64'd9763909481373, - 64'd152465666597786, - 64'd4973942635102, - 64'd152787603191753, - 64'd729699476620, - 64'd151191882518354, 64'd2985818768773, - 64'd147941048171172, 64'd6193952317251, - 64'd143284714725683, 64'd8919570676754, - 64'd137458139359128, 64'd11190320031248, - 64'd130681150796010, 64'd13035931862094, - 64'd123157403467911, 64'd14487593541614, - 64'd115073924849368, 64'd15577380779578, - 64'd106600924388957, 64'd16337751058586, - 64'd97891833242094, 64'd16801096554637},
		'{- 64'd16661173520135, - 64'd67604904587707, - 64'd46932306946327, - 64'd58666327761395, - 64'd72791968326060, - 64'd50139480307340, - 64'd94481366958141, - 64'd42076947065871, - 64'd112262382465842, - 64'd34518947358519, - 64'd126411729164527, - 64'd27494407471536, - 64'd137215677493413, - 64'd21022035995946, - 64'd144965326781880, - 64'd15111388452564, - 64'd149952417573864, - 64'd9763909481373, - 64'd152465666597786, - 64'd4973942635102, - 64'd152787603191753, - 64'd729699476620, - 64'd151191882518354, 64'd2985818768773, - 64'd147941048171172, 64'd6193952317251, - 64'd143284714725683, 64'd8919570676754, - 64'd137458139359128, 64'd11190320031248, - 64'd130681150796010, 64'd13035931862094, - 64'd123157403467911, 64'd14487593541614, - 64'd115073924849368, 64'd15577380779578, - 64'd106600924388957, 64'd16337751058586, - 64'd97891833242094, 64'd16801096554637}};
	localparam logic signed[63:0] Ffi[0:1][0:39] = '{
		'{64'd363978915924475, - 64'd49115498086959, 64'd337249040609096, - 64'd51540235037469, 64'd309762650084378, - 64'd53024660207131, 64'd281953232772926, - 64'd53669663522991, 64'd254203328051453, - 64'd53573665130579, 64'd226846281624461, - 64'd52831719270158, 64'd200168382820128, - 64'd51534773027261, 64'd174411309169022, - 64'd49769069442666, 64'd149774809307364, - 64'd47615684025719, 64'd126419561055001, - 64'd45150183464151, 64'd104470147366645, - 64'd42442395242206, 64'd84018098666250, - 64'd39556276946533, 64'd65124955782048, - 64'd36549874236225, 64'd47825313246755, - 64'd33475356760732, 64'd32129808065913, - 64'd30379121709495, 64'd18028024148230, - 64'd27301955153229, 64'd5491287403838, - 64'd24279241873493, - 64'd5524668974162, - 64'd21341214960134, - 64'd15077185339646, - 64'd18513237072459, - 64'd23234314970514, - 64'd15816105897687},
		'{- 64'd363978915924475, 64'd49115498086959, - 64'd337249040609096, 64'd51540235037469, - 64'd309762650084377, 64'd53024660207131, - 64'd281953232772926, 64'd53669663522991, - 64'd254203328051453, 64'd53573665130579, - 64'd226846281624461, 64'd52831719270158, - 64'd200168382820128, 64'd51534773027261, - 64'd174411309169022, 64'd49769069442666, - 64'd149774809307364, 64'd47615684025719, - 64'd126419561055001, 64'd45150183464151, - 64'd104470147366645, 64'd42442395242206, - 64'd84018098666250, 64'd39556276946533, - 64'd65124955782048, 64'd36549874236225, - 64'd47825313246755, 64'd33475356760732, - 64'd32129808065913, 64'd30379121709495, - 64'd18028024148230, 64'd27301955153229, - 64'd5491287403838, 64'd24279241873493, 64'd5524668974162, 64'd21341214960134, 64'd15077185339647, 64'd18513237072459, 64'd23234314970514, 64'd15816105897687}};
	localparam logic signed[63:0] Fbr[0:1][0:39] = '{
		'{- 64'd16661173520135, 64'd67604904587707, - 64'd46932306946327, 64'd58666327761395, - 64'd72791968326060, 64'd50139480307340, - 64'd94481366958141, 64'd42076947065871, - 64'd112262382465842, 64'd34518947358519, - 64'd126411729164527, 64'd27494407471536, - 64'd137215677493413, 64'd21022035995946, - 64'd144965326781880, 64'd15111388452564, - 64'd149952417573864, 64'd9763909481373, - 64'd152465666597786, 64'd4973942635102, - 64'd152787603191753, 64'd729699476620, - 64'd151191882518354, - 64'd2985818768773, - 64'd147941048171172, - 64'd6193952317251, - 64'd143284714725683, - 64'd8919570676754, - 64'd137458139359128, - 64'd11190320031248, - 64'd130681150796010, - 64'd13035931862094, - 64'd123157403467911, - 64'd14487593541614, - 64'd115073924849368, - 64'd15577380779578, - 64'd106600924388957, - 64'd16337751058586, - 64'd97891833242094, - 64'd16801096554637},
		'{- 64'd16661173520135, 64'd67604904587707, - 64'd46932306946327, 64'd58666327761395, - 64'd72791968326060, 64'd50139480307340, - 64'd94481366958141, 64'd42076947065871, - 64'd112262382465842, 64'd34518947358519, - 64'd126411729164527, 64'd27494407471536, - 64'd137215677493413, 64'd21022035995946, - 64'd144965326781880, 64'd15111388452564, - 64'd149952417573864, 64'd9763909481373, - 64'd152465666597786, 64'd4973942635102, - 64'd152787603191753, 64'd729699476620, - 64'd151191882518354, - 64'd2985818768773, - 64'd147941048171172, - 64'd6193952317251, - 64'd143284714725683, - 64'd8919570676754, - 64'd137458139359128, - 64'd11190320031248, - 64'd130681150796010, - 64'd13035931862094, - 64'd123157403467911, - 64'd14487593541614, - 64'd115073924849368, - 64'd15577380779578, - 64'd106600924388957, - 64'd16337751058586, - 64'd97891833242094, - 64'd16801096554637}};
	localparam logic signed[63:0] Fbi[0:1][0:39] = '{
		'{64'd363978915924475, 64'd49115498086959, 64'd337249040609096, 64'd51540235037469, 64'd309762650084378, 64'd53024660207131, 64'd281953232772926, 64'd53669663522991, 64'd254203328051453, 64'd53573665130579, 64'd226846281624461, 64'd52831719270158, 64'd200168382820128, 64'd51534773027261, 64'd174411309169022, 64'd49769069442666, 64'd149774809307364, 64'd47615684025719, 64'd126419561055001, 64'd45150183464151, 64'd104470147366645, 64'd42442395242206, 64'd84018098666250, 64'd39556276946533, 64'd65124955782048, 64'd36549874236225, 64'd47825313246755, 64'd33475356760732, 64'd32129808065913, 64'd30379121709495, 64'd18028024148230, 64'd27301955153229, 64'd5491287403838, 64'd24279241873493, - 64'd5524668974162, 64'd21341214960134, - 64'd15077185339646, 64'd18513237072459, - 64'd23234314970514, 64'd15816105897687},
		'{- 64'd363978915924475, - 64'd49115498086959, - 64'd337249040609096, - 64'd51540235037469, - 64'd309762650084377, - 64'd53024660207131, - 64'd281953232772926, - 64'd53669663522991, - 64'd254203328051453, - 64'd53573665130579, - 64'd226846281624461, - 64'd52831719270158, - 64'd200168382820128, - 64'd51534773027261, - 64'd174411309169022, - 64'd49769069442666, - 64'd149774809307364, - 64'd47615684025719, - 64'd126419561055001, - 64'd45150183464151, - 64'd104470147366645, - 64'd42442395242206, - 64'd84018098666250, - 64'd39556276946533, - 64'd65124955782048, - 64'd36549874236225, - 64'd47825313246755, - 64'd33475356760732, - 64'd32129808065913, - 64'd30379121709495, - 64'd18028024148230, - 64'd27301955153229, - 64'd5491287403838, - 64'd24279241873493, 64'd5524668974162, - 64'd21341214960134, 64'd15077185339647, - 64'd18513237072459, 64'd23234314970514, - 64'd15816105897687}};
	localparam logic signed[63:0] hf[0:599] = {64'd12785266196480, - 64'd156027043840, 64'd12553857007616, - 64'd439507386368, 64'd12197550882816, - 64'd681675587584, 64'd11736547590144, - 64'd884790525952, 64'd11189771829248, - 64'd1051304525824, 64'd10574809268224, - 64'd1183809011712, 64'd9907850969088, - 64'd1284984930304, 64'd9203676610560, - 64'd1357558054912, 64'd8475652390912, - 64'd1404260712448, 64'd7735742562304, - 64'd1427796656128, 64'd6994541936640, - 64'd1430811443200, 64'd6261319401472, - 64'd1415868055552, 64'd5544070873088, - 64'd1385424879616, 64'd4849583783936, - 64'd1341819715584, 64'd4183505764352, - 64'd1287255490560, 64'd3550419877888, - 64'd1223790952448, 64'd2953923526656, - 64'd1153333198848, 64'd2396708405248, - 64'd1077633810432, 64'd1880643600384, - 64'd998286622720, 64'd1406855020544, - 64'd916728512512, 64'd975806988288, - 64'd834241495040, 64'd587379965952, - 64'd751956459520, 64'd240945954816, - 64'd670858674176, - 64'd64559341568, - 64'd591793881088, - 64'd330568138752, - 64'd515475865600, - 64'd558816428032, - 64'd442494124032, - 64'd751284125696, - 64'd373322481664, - 64'd910139850752, - 64'd308328005632, - 64'd1037690339328, - 64'd247779901440, - 64'd1136334733312, - 64'd191858655232, - 64'd1208523161600, - 64'd140665044992, - 64'd1256720564224, - 64'd94229028864, - 64'd1283374317568, - 64'd52518301696, - 64'd1290886053888, - 64'd15446620160, - 64'd1281588723712, 64'd17118325760, - 64'd1257726017536, 64'd45347446784, - 64'd1221436112896, 64'd69443256320, - 64'd1174739353600, 64'd89633398784, - 64'd1119527763968, 64'd106164649984, - 64'd1057558233088, 64'd119297458176, - 64'd990448123904, 64'd129301045248, - 64'd919673176064, 64'd136448958464, - 64'd846566981632, 64'd141015154688, - 64'd772322951168, 64'd143270625280, - 64'd697997328384, 64'd143480389632, - 64'd624513384448, 64'd141901037568, - 64'd552667250688, 64'd138778640384, - 64'd483134013440, 64'd134347014144, - 64'd416474759168, 64'd128826466304, - 64'd353144307712, 64'd122422779904, - 64'd293498847232, 64'd115326484480, - 64'd237804290048, 64'd107712503808, - 64'd186244251648, 64'd99739951104, - 64'd138928324608, 64'd91552186368, - 64'd95900065792, 64'd83277062144, - 64'd57144852480, 64'd75027292160, - 64'd22597429248, 64'd66901004288, 64'd7850891264, 64'd58982383616, 64'd34345375744, 64'd51342397440, 64'd57061462016, 64'd44039593984, 64'd76198764544, 64'd37120970752, 64'd91975589888, 64'd30622838784, 64'd104623857664, 64'd24571756544, 64'd114384543744, 64'd18985422848, 64'd121503555584, 64'd13873581056, 64'd126228111360, 64'd9238916096, 64'd128803520512, 64'd5077907456, 64'd129470414848, 64'd1381665152, 64'd128462381056, - 64'd1863285376, 64'd126003994624, - 64'd4674255360, 64'd122309197824, - 64'd7071693312, 64'd117580013568, - 64'd9078538240, 64'd112005570560, - 64'd10719621120, 64'd105761439744, - 64'd12021117952, 64'd99009167360, - 64'd13010063360, 64'd91896070144, - 64'd13713903616, 64'd84555235328, - 64'd14160113664, 64'd77105692672, - 64'd14375848960, 64'd69652725760, - 64'd14387657728, 64'd62288318464, - 64'd14221230080, 64'd55091728384, - 64'd13901189120, 64'd48130088960, - 64'd13450929152, 64'd41459154944, - 64'd12892477440, 64'd35124047872, - 64'd12246400000, 64'd29160044544, - 64'd11531735040, 64'd23593392128, - 64'd10765949952, 64'd18442135552, - 64'd9964929024, 64'd13716925440, - 64'd9142975488, 64'd9421835264, - 64'd8312838656, 64'd5555136512, - 64'd7485752320, 64'd2110055680, - 64'd6671490048, - 64'd924499968, - 64'd5878430208, - 64'd3563261440, - 64'd5113628672, - 64'd5823955456, - 64'd4382900736, - 64'd7726706688, - 64'd3690905344, - 64'd9293489152, - 64'd3041236992, - 64'd10547617792, - 64'd2436513536, - 64'd11513296896, - 64'd1878470016, - 64'd12215205888, - 64'd1368047616, - 64'd12678137856, - 64'd905483520, - 64'd12926682112, - 64'd490396960, - 64'd12984944640, - 64'd121872168, - 64'd12876317696, 64'd201462592, - 64'd12623277056, 64'd481360352, - 64'd12247225344, 64'd719885696, - 64'd11768368128, 64'd919349888, - 64'd11205610496, 64'd1082251136, - 64'd10576494592, 64'd1211220480, - 64'd9897156608, 64'd1308972160, - 64'd9182302208, 64'd1378260480, - 64'd8445213184, 64'd1421840000, - 64'd7697760768, 64'd1442432384, - 64'd6950439936, 64'd1442696960, - 64'd6212413952, 64'd1425205632, - 64'd5491571712, 64'd1392422656, - 64'd4794590720, 64'd1346688128, - 64'd4127010304, 64'd1290204544, - 64'd3493306368, 64'd1225027584, - 64'd2896971776, 64'd1153059200, - 64'd2340597760, 64'd1076043776, - 64'd1825956736, 64'd995566912, - 64'd1354083200, 64'd913055616, - 64'd925356032, 64'd829781248, - 64'd539575552, 64'd746863424, - 64'd196040048, 64'd665275584, 64'd106382320, 64'd585851456, 64'd369184992, 64'd509292608, 64'd594158976, 64'd436176448, 64'd783332992, 64'd366965088, 64'd938918592, 64'd302013984, 64'd1063259776, 64'd241581328, 64'd1158787200, 64'd185837040, 64'd1227977856, 64'd134871952, 64'd1273318400, 64'd88706664, 64'd1297273088, 64'd47300204, 64'd1302257152, 64'd10558347, 64'd1290612480, - 64'd21658510, 64'd1264589056, - 64'd49527868, 64'd1226327936, - 64'd73258144, 64'd1177849600, - 64'd93082192, 64'd1121043840, - 64'd109251360, 64'd1057663488, - 64'd122030048, 64'd989320000, - 64'd131690800, 64'd917481792, - 64'd138509952, 64'd843473920, - 64'd142763728, 64'd768480512, - 64'd144724880, 64'd693547584, - 64'd144659744, 64'd619587968, - 64'd142825824, 64'd547386944, - 64'd139469744, 64'd477608608, - 64'd134825568, 64'd410803200, - 64'd129113520, 64'd347414752, - 64'd122539048, 64'd287789056, - 64'd115292192, 64'd232181904, - 64'd107547136, 64'd180767248, - 64'd99462152, 64'd133645568, - 64'd91179608, 64'd90851840, - 64'd82826288, 64'd52363464, - 64'd74513760, 64'd18107806, - 64'd66338984, - 64'd12030560, - 64'd58384920, - 64'd38203012, - 64'd50721320, - 64'd60590476, - 64'd43405520, - 64'd79397440, - 64'd36483336, - 64'd94846480, - 64'd29989930, - 64'd107173224, - 64'd23950750, - 64'd116621800, - 64'd18382436, - 64'd123440760, - 64'd13293740, - 64'd127879480, - 64'd8686411, - 64'd130184976, - 64'd4556064, - 64'd130599184, - 64'd893008, - 64'd129356608, 64'd2316958, - 64'd126682408, 64'd5091802, - 64'd122790808, 64'd7452562, - 64'd117883832, 64'd9422696, - 64'd112150392, 64'd11027491, - 64'd105765632, 64'd12293516, - 64'd98890488, 64'd13248137, - 64'd91671544, 64'd13919077, - 64'd84241032, 64'd14334034, - 64'd76717032, 64'd14520339, - 64'd69203816, 64'd14504671, - 64'd61792308, 64'd14312810, - 64'd54560672, 64'd13969434, - 64'd47574952, 64'd13497956, - 64'd40889812, 64'd12920396, - 64'd34549288, 64'd12257289, - 64'd28587616, 64'd11527617, - 64'd23030032, 64'd10748778, - 64'd17893614, 64'd9936567, - 64'd13188102, 64'd9105190, - 64'd8916710, 64'd8267287, - 64'd5076912, 64'd7433978, - 64'd1661199, 64'd6614918, 64'd1342196, 64'd5818363, 64'd3948613, 64'd5051247, 64'd6176326, 64'd4319264, 64'd8045947, 64'd3626954, 64'd9579874, 64'd2977797, 64'd10801792, 64'd2374299, 64'd11736218, 64'd1818090, 64'd12408095, 64'd1310012, 64'd12842430, 64'd850207, 64'd13063983, 64'd438210, 64'd13096987, 64'd73024, 64'd12964924, - 64'd246794, 64'd12690328, - 64'd523065, 64'd12294629, - 64'd757910, 64'd11798031, - 64'd953693, 64'd11219415, - 64'd1112958, 64'd10576281, - 64'd1238374, 64'd9884702, - 64'd1332689, 64'd9159312, - 64'd1398685, 64'd8413304, - 64'd1439138, 64'd7658454, - 64'd1456788, 64'd6905156, - 64'd1454306, 64'd6162466, - 64'd1434274, 64'd5438165, - 64'd1399160, 64'd4738819, - 64'd1351308, 64'd4069858, - 64'd1292918, 64'd3435651, - 64'd1226043, 64'd2839585, - 64'd1152579, 64'd2284151, - 64'd1074263, 64'd1771024, - 64'd992673, 64'd1301147, - 64'd909224, 64'd874814, - 64'd825179, 64'd491746, - 64'd741644, 64'd151166, - 64'd659582, - 64'd148124, - 64'd579813, - 64'd407678, - 64'd503027, - 64'd629342, - 64'd429790, - 64'd815194, - 64'd360551, - 64'd967486, - 64'd295655, - 64'd1088600, - 64'd235349, - 64'd1180998, - 64'd179791, - 64'd1247183, - 64'd129063, - 64'd1289663, - 64'd83177, - 64'd1310918, - 64'd42081, - 64'd1313378, - 64'd5675, - 64'd1299391, 64'd26188, - 64'd1271215, 64'd53693, - 64'd1230992, 64'd77054, - 64'd1180744, 64'd96509, - 64'd1122356, 64'd112314, - 64'd1057579, 64'd124737, - 64'd988016, 64'd134053, - 64'd915129, 64'd140543, - 64'd840234, 64'd144484, - 64'd764506, 64'd146151, - 64'd688980, 64'd145811, - 64'd614559, 64'd143724, - 64'd542016, 64'd140135, - 64'd472006, 64'd135279, - 64'd405066, 64'd129377, - 64'd341631, 64'd122633, - 64'd282036, 64'd115237, - 64'd226526, 64'd107363, - 64'd175266, 64'd99167, - 64'd128347, 64'd90791, - 64'd85795, 64'd82361, - 64'd47580, 64'd73988, - 64'd13622, 64'd65766, 64'd16202, 64'd57778, 64'd42048, 64'd50092, 64'd64103, 64'd42765, 64'd82577, 64'd35840, 64'd97696, 64'd29353, 64'd109700, 64'd23326, 64'd118835, 64'd17777, 64'd125353, 64'd12712, 64'd129505, 64'd8133, 64'd131541, 64'd4034, 64'd131703, 64'd405, 64'd130226, - 64'd2770, 64'd127337, - 64'd5508, 64'd123250, - 64'd7832, 64'd118166, - 64'd9765, 64'd112275, - 64'd11333, 64'd105751, - 64'd12563, 64'd98754, - 64'd13483, 64'd91431, - 64'd14121, 64'd83912, - 64'd14505, 64'd76315, - 64'd14662, 64'd68743, - 64'd14619, 64'd61286, - 64'd14402, 64'd54021, - 64'd14035, 64'd47012, - 64'd13542, 64'd40314, - 64'd12946, 64'd33969, - 64'd12266, 64'd28011, - 64'd11521, 64'd22463, - 64'd10730, 64'd17343, - 64'd9906, 64'd12658, - 64'd9066, 64'd8411, - 64'd8220, 64'd4598, - 64'd7381, 64'd1213, - 64'd6557, - 64'd1759, - 64'd5757, - 64'd4333, - 64'd4988, - 64'd6527, - 64'd4255, - 64'd8363, - 64'd3562, - 64'd9864, - 64'd2914};
	localparam logic signed[63:0] hb[0:599] = {64'd12785266196480, 64'd156027043840, 64'd12553857007616, 64'd439507386368, 64'd12197550882816, 64'd681675587584, 64'd11736547590144, 64'd884790525952, 64'd11189771829248, 64'd1051304525824, 64'd10574809268224, 64'd1183809011712, 64'd9907850969088, 64'd1284984930304, 64'd9203676610560, 64'd1357558054912, 64'd8475652390912, 64'd1404260712448, 64'd7735742562304, 64'd1427796656128, 64'd6994541936640, 64'd1430811443200, 64'd6261319401472, 64'd1415868055552, 64'd5544070873088, 64'd1385424879616, 64'd4849583783936, 64'd1341819715584, 64'd4183505764352, 64'd1287255490560, 64'd3550419877888, 64'd1223790952448, 64'd2953923526656, 64'd1153333198848, 64'd2396708405248, 64'd1077633810432, 64'd1880643600384, 64'd998286622720, 64'd1406855020544, 64'd916728512512, 64'd975806988288, 64'd834241495040, 64'd587379965952, 64'd751956459520, 64'd240945954816, 64'd670858674176, - 64'd64559341568, 64'd591793881088, - 64'd330568138752, 64'd515475865600, - 64'd558816428032, 64'd442494124032, - 64'd751284125696, 64'd373322481664, - 64'd910139850752, 64'd308328005632, - 64'd1037690339328, 64'd247779901440, - 64'd1136334733312, 64'd191858655232, - 64'd1208523161600, 64'd140665044992, - 64'd1256720564224, 64'd94229028864, - 64'd1283374317568, 64'd52518301696, - 64'd1290886053888, 64'd15446620160, - 64'd1281588723712, - 64'd17118325760, - 64'd1257726017536, - 64'd45347446784, - 64'd1221436112896, - 64'd69443256320, - 64'd1174739353600, - 64'd89633398784, - 64'd1119527763968, - 64'd106164649984, - 64'd1057558233088, - 64'd119297458176, - 64'd990448123904, - 64'd129301045248, - 64'd919673176064, - 64'd136448958464, - 64'd846566981632, - 64'd141015154688, - 64'd772322951168, - 64'd143270625280, - 64'd697997328384, - 64'd143480389632, - 64'd624513384448, - 64'd141901037568, - 64'd552667250688, - 64'd138778640384, - 64'd483134013440, - 64'd134347014144, - 64'd416474759168, - 64'd128826466304, - 64'd353144307712, - 64'd122422779904, - 64'd293498847232, - 64'd115326484480, - 64'd237804290048, - 64'd107712503808, - 64'd186244251648, - 64'd99739951104, - 64'd138928324608, - 64'd91552186368, - 64'd95900065792, - 64'd83277062144, - 64'd57144852480, - 64'd75027292160, - 64'd22597429248, - 64'd66901004288, 64'd7850891264, - 64'd58982383616, 64'd34345375744, - 64'd51342397440, 64'd57061462016, - 64'd44039593984, 64'd76198764544, - 64'd37120970752, 64'd91975589888, - 64'd30622838784, 64'd104623857664, - 64'd24571756544, 64'd114384543744, - 64'd18985422848, 64'd121503555584, - 64'd13873581056, 64'd126228111360, - 64'd9238916096, 64'd128803520512, - 64'd5077907456, 64'd129470414848, - 64'd1381665152, 64'd128462381056, 64'd1863285376, 64'd126003994624, 64'd4674255360, 64'd122309197824, 64'd7071693312, 64'd117580013568, 64'd9078538240, 64'd112005570560, 64'd10719621120, 64'd105761439744, 64'd12021117952, 64'd99009167360, 64'd13010063360, 64'd91896070144, 64'd13713903616, 64'd84555235328, 64'd14160113664, 64'd77105692672, 64'd14375848960, 64'd69652725760, 64'd14387657728, 64'd62288318464, 64'd14221230080, 64'd55091728384, 64'd13901189120, 64'd48130088960, 64'd13450929152, 64'd41459154944, 64'd12892477440, 64'd35124047872, 64'd12246400000, 64'd29160044544, 64'd11531735040, 64'd23593392128, 64'd10765949952, 64'd18442135552, 64'd9964929024, 64'd13716925440, 64'd9142975488, 64'd9421835264, 64'd8312838656, 64'd5555136512, 64'd7485752320, 64'd2110055680, 64'd6671490048, - 64'd924499968, 64'd5878430208, - 64'd3563261440, 64'd5113628672, - 64'd5823955456, 64'd4382900736, - 64'd7726706688, 64'd3690905344, - 64'd9293489152, 64'd3041236992, - 64'd10547617792, 64'd2436513536, - 64'd11513296896, 64'd1878470016, - 64'd12215205888, 64'd1368047616, - 64'd12678137856, 64'd905483520, - 64'd12926682112, 64'd490396960, - 64'd12984944640, 64'd121872168, - 64'd12876317696, - 64'd201462592, - 64'd12623277056, - 64'd481360352, - 64'd12247225344, - 64'd719885696, - 64'd11768368128, - 64'd919349888, - 64'd11205610496, - 64'd1082251136, - 64'd10576494592, - 64'd1211220480, - 64'd9897156608, - 64'd1308972160, - 64'd9182302208, - 64'd1378260480, - 64'd8445213184, - 64'd1421840000, - 64'd7697760768, - 64'd1442432384, - 64'd6950439936, - 64'd1442696960, - 64'd6212413952, - 64'd1425205632, - 64'd5491571712, - 64'd1392422656, - 64'd4794590720, - 64'd1346688128, - 64'd4127010304, - 64'd1290204544, - 64'd3493306368, - 64'd1225027584, - 64'd2896971776, - 64'd1153059200, - 64'd2340597760, - 64'd1076043776, - 64'd1825956736, - 64'd995566912, - 64'd1354083200, - 64'd913055616, - 64'd925356032, - 64'd829781248, - 64'd539575552, - 64'd746863424, - 64'd196040048, - 64'd665275584, 64'd106382320, - 64'd585851456, 64'd369184992, - 64'd509292608, 64'd594158976, - 64'd436176448, 64'd783332992, - 64'd366965088, 64'd938918592, - 64'd302013984, 64'd1063259776, - 64'd241581328, 64'd1158787200, - 64'd185837040, 64'd1227977856, - 64'd134871952, 64'd1273318400, - 64'd88706664, 64'd1297273088, - 64'd47300204, 64'd1302257152, - 64'd10558347, 64'd1290612480, 64'd21658510, 64'd1264589056, 64'd49527868, 64'd1226327936, 64'd73258144, 64'd1177849600, 64'd93082192, 64'd1121043840, 64'd109251360, 64'd1057663488, 64'd122030048, 64'd989320000, 64'd131690800, 64'd917481792, 64'd138509952, 64'd843473920, 64'd142763728, 64'd768480512, 64'd144724880, 64'd693547584, 64'd144659744, 64'd619587968, 64'd142825824, 64'd547386944, 64'd139469744, 64'd477608608, 64'd134825568, 64'd410803200, 64'd129113520, 64'd347414752, 64'd122539048, 64'd287789056, 64'd115292192, 64'd232181904, 64'd107547136, 64'd180767248, 64'd99462152, 64'd133645568, 64'd91179608, 64'd90851840, 64'd82826288, 64'd52363464, 64'd74513760, 64'd18107806, 64'd66338984, - 64'd12030560, 64'd58384920, - 64'd38203012, 64'd50721320, - 64'd60590476, 64'd43405520, - 64'd79397440, 64'd36483336, - 64'd94846480, 64'd29989930, - 64'd107173224, 64'd23950750, - 64'd116621800, 64'd18382436, - 64'd123440760, 64'd13293740, - 64'd127879480, 64'd8686411, - 64'd130184976, 64'd4556064, - 64'd130599184, 64'd893008, - 64'd129356608, - 64'd2316958, - 64'd126682408, - 64'd5091802, - 64'd122790808, - 64'd7452562, - 64'd117883832, - 64'd9422696, - 64'd112150392, - 64'd11027491, - 64'd105765632, - 64'd12293516, - 64'd98890488, - 64'd13248137, - 64'd91671544, - 64'd13919077, - 64'd84241032, - 64'd14334034, - 64'd76717032, - 64'd14520339, - 64'd69203816, - 64'd14504671, - 64'd61792308, - 64'd14312810, - 64'd54560672, - 64'd13969434, - 64'd47574952, - 64'd13497956, - 64'd40889812, - 64'd12920396, - 64'd34549288, - 64'd12257289, - 64'd28587616, - 64'd11527617, - 64'd23030032, - 64'd10748778, - 64'd17893614, - 64'd9936567, - 64'd13188102, - 64'd9105190, - 64'd8916710, - 64'd8267287, - 64'd5076912, - 64'd7433978, - 64'd1661199, - 64'd6614918, 64'd1342196, - 64'd5818363, 64'd3948613, - 64'd5051247, 64'd6176326, - 64'd4319264, 64'd8045947, - 64'd3626954, 64'd9579874, - 64'd2977797, 64'd10801792, - 64'd2374299, 64'd11736218, - 64'd1818090, 64'd12408095, - 64'd1310012, 64'd12842430, - 64'd850207, 64'd13063983, - 64'd438210, 64'd13096987, - 64'd73024, 64'd12964924, 64'd246794, 64'd12690328, 64'd523065, 64'd12294629, 64'd757910, 64'd11798031, 64'd953693, 64'd11219415, 64'd1112958, 64'd10576281, 64'd1238374, 64'd9884702, 64'd1332689, 64'd9159312, 64'd1398685, 64'd8413304, 64'd1439138, 64'd7658454, 64'd1456788, 64'd6905156, 64'd1454306, 64'd6162466, 64'd1434274, 64'd5438165, 64'd1399160, 64'd4738819, 64'd1351308, 64'd4069858, 64'd1292918, 64'd3435651, 64'd1226043, 64'd2839585, 64'd1152579, 64'd2284151, 64'd1074263, 64'd1771024, 64'd992673, 64'd1301147, 64'd909224, 64'd874814, 64'd825179, 64'd491746, 64'd741644, 64'd151166, 64'd659582, - 64'd148124, 64'd579813, - 64'd407678, 64'd503027, - 64'd629342, 64'd429790, - 64'd815194, 64'd360551, - 64'd967486, 64'd295655, - 64'd1088600, 64'd235349, - 64'd1180998, 64'd179791, - 64'd1247183, 64'd129063, - 64'd1289663, 64'd83177, - 64'd1310918, 64'd42081, - 64'd1313378, 64'd5675, - 64'd1299391, - 64'd26188, - 64'd1271215, - 64'd53693, - 64'd1230992, - 64'd77054, - 64'd1180744, - 64'd96509, - 64'd1122356, - 64'd112314, - 64'd1057579, - 64'd124737, - 64'd988016, - 64'd134053, - 64'd915129, - 64'd140543, - 64'd840234, - 64'd144484, - 64'd764506, - 64'd146151, - 64'd688980, - 64'd145811, - 64'd614559, - 64'd143724, - 64'd542016, - 64'd140135, - 64'd472006, - 64'd135279, - 64'd405066, - 64'd129377, - 64'd341631, - 64'd122633, - 64'd282036, - 64'd115237, - 64'd226526, - 64'd107363, - 64'd175266, - 64'd99167, - 64'd128347, - 64'd90791, - 64'd85795, - 64'd82361, - 64'd47580, - 64'd73988, - 64'd13622, - 64'd65766, 64'd16202, - 64'd57778, 64'd42048, - 64'd50092, 64'd64103, - 64'd42765, 64'd82577, - 64'd35840, 64'd97696, - 64'd29353, 64'd109700, - 64'd23326, 64'd118835, - 64'd17777, 64'd125353, - 64'd12712, 64'd129505, - 64'd8133, 64'd131541, - 64'd4034, 64'd131703, - 64'd405, 64'd130226, 64'd2770, 64'd127337, 64'd5508, 64'd123250, 64'd7832, 64'd118166, 64'd9765, 64'd112275, 64'd11333, 64'd105751, 64'd12563, 64'd98754, 64'd13483, 64'd91431, 64'd14121, 64'd83912, 64'd14505, 64'd76315, 64'd14662, 64'd68743, 64'd14619, 64'd61286, 64'd14402, 64'd54021, 64'd14035, 64'd47012, 64'd13542, 64'd40314, 64'd12946, 64'd33969, 64'd12266, 64'd28011, 64'd11521, 64'd22463, 64'd10730, 64'd17343, 64'd9906, 64'd12658, 64'd9066, 64'd8411, 64'd8220, 64'd4598, 64'd7381, 64'd1213, 64'd6557, - 64'd1759, 64'd5757, - 64'd4333, 64'd4988, - 64'd6527, 64'd4255, - 64'd8363, 64'd3562, - 64'd9864, 64'd2914};
endpackage
`endif
